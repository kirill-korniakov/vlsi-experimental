# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2008, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use.  This file contains valuable trade secrets and    *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *          NGLibraryCreator Development_version build 200801281737           *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on server08.nangate.com for user Paulo Butzen (pbu).
# Local time is now Fri, 22 Feb 2008, 21:19:06.
# Main process id is 11136.

VERSION 5.3 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

# Export LEF: 6 routing layers requested in librarytemplate, but only 3 metal layer(s) available.
LAYER M1
  TYPE ROUTING ;
  WIDTH 0.065 ;
  SPACING 0.065 ;
  PITCH 0.14 ;
  DIRECTION HORIZONTAL ;
  RESISTANCE RPERSQ 0.38 ;
  THICKNESS 0.13 ;
  CAPACITANCE CPERSQDIST 0.001 ;
  EDGECAPACITANCE 5.00e-04 ;
END M1

LAYER V1
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.065 ;
END V1

LAYER M2
  TYPE ROUTING ;
  WIDTH 0.07 ;
  SPACING 0.07 ;
  PITCH 0.19 ;
  DIRECTION VERTICAL ;
  RESISTANCE RPERSQ 0.25 ;
  THICKNESS 0.14 ;
  CAPACITANCE CPERSQDIST 0.001 ;
  EDGECAPACITANCE 5.00e-04 ;
END M2

LAYER V2
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.065 ;
END V2

LAYER M3
  TYPE ROUTING ;
  WIDTH 0.07 ;
  SPACING 0.07 ;
  PITCH 0.14 ;
  DIRECTION HORIZONTAL ;
  RESISTANCE RPERSQ 0.25 ;
  THICKNESS 0.14 ;
  CAPACITANCE CPERSQDIST 0.001 ;
  EDGECAPACITANCE 5.00e-04 ;
END M3

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA Via1 DEFAULT
  RESISTANCE 1 ;
  LAYER V1 ;
    RECT -0.03 -0.03 0.035 0.035 ;
  LAYER M1 ;
    RECT -0.065 -0.065 0.07 0.07 ;
  LAYER M2 ;
    RECT -0.065 -0.065 0.07 0.07 ;
END Via1

VIA Via2 DEFAULT
  RESISTANCE 1 ;
  LAYER V2 ;
    RECT -0.03 -0.03 0.035 0.035 ;
  LAYER M2 ;
    RECT -0.065 -0.065 0.07 0.07 ;
  LAYER M3 ;
    RECT -0.065 -0.065 0.07 0.07 ;
END Via2

VIARULE Via1Array GENERATE
  LAYER M1 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER M2 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER V1 ;
    RECT -0.03 -0.03 0.035 0.035 ;
    SPACING 0.14 BY 0.14 ;
END Via1Array

VIARULE Via2Array GENERATE
  LAYER M2 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER M3 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER V2 ;
    RECT -0.03 -0.03 0.035 0.035 ;
    SPACING 0.14 BY 0.14 ;
END Via2Array

VIARULE TURNM1 GENERATE
  LAYER M1 ;
    DIRECTION vertical ;
  LAYER M1 ;
    DIRECTION horizontal ;
END TURNM1

VIARULE TURNM2 GENERATE
  LAYER M2 ;
    DIRECTION vertical ;
  LAYER M2 ;
    DIRECTION horizontal ;
END TURNM2

VIARULE TURNM3 GENERATE
  LAYER M3 ;
    DIRECTION vertical ;
  LAYER M3 ;
    DIRECTION horizontal ;
END TURNM3

SPACING
  SAMENET M1 M1 0.065 ;
  SAMENET M2 M2 0.07 ;
  SAMENET M3 M3 0.07 ;
  SAMENET V1 V1 0.075 ;
  SAMENET V2 V2 0.075 ;
  SAMENET V1 V2 0.0 STACK ;
END SPACING

SITE Free_OMC_Si2_PDK45nm
  SYMMETRY y ;
  CLASS core ;
  SIZE 0.19 BY 1.4 ;
END Free_OMC_Si2_PDK45nm

MACRO XNOR2_X1
  CLASS core ;
  FOREIGN XNOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.9 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.205 0.57 0.695 0.57 0.695 0.5 0.76 0.5 0.76 0.635 0.27 0.635 0.27 0.705 0.205 0.705  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.31 1.315 0.31 1.125 0.375 1.125 0.375 1.315 1.41 1.315 1.41 1.125 1.475 1.125 1.475 1.315 1.9 1.315 1.9 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.9 -0.085 1.9 0.085 1.575 0.085 1.575 0.15 1.51 0.15 1.51 0.365 1.445 0.365 1.445 0.085 0.3 0.085 0.3 0.33 0.235 0.33 0.235 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.355 0.37 0.49 0.37 0.49 0.505 0.355 0.505  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.58 0.245 1.73 0.245 1.73 1.155 1.58 1.155  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.555 0.86 0.62 0.86 0.62 1.155 0.555 1.155  ;
        POLYGON 0.05 0.21 0.115 0.21 0.115 0.77 0.33 0.77 0.33 0.73 0.855 0.73 0.855 0.475 0.92 0.475 0.92 0.795 0.78 0.795 0.78 0.995 0.715 0.995 0.715 0.795 0.39 0.795 0.39 0.835 0.19 0.835 0.19 1.155 0.05 1.155  ;
        POLYGON 1.08 1.055 1.115 1.055 1.115 0.345 1.115 0.28 1.25 0.28 1.25 0.345 1.215 0.345 1.215 0.38 1.18 0.38 1.18 1.055 1.215 1.055 1.215 1.12 1.08 1.12  ;
        POLYGON 0.555 0.15 1.38 0.15 1.38 0.54 1.315 0.54 1.315 0.215 0.62 0.215 0.62 0.505 0.555 0.505  ;
        POLYGON 0.98 1.055 1.015 1.055 1.015 1.185 1.28 1.185 1.28 0.93 1.45 0.93 1.45 0.86 1.515 0.86 1.515 0.995 1.345 0.995 1.345 1.25 0.95 1.25 0.95 1.155 0.915 1.155 0.915 0.86 0.985 0.86 0.985 0.41 0.85 0.41 0.85 0.345 0.815 0.345 0.815 0.28 0.95 0.28 0.95 0.345 1.05 0.345 1.05 0.925 0.98 0.925  ;
  END
END XNOR2_X1

MACRO XNOR2_X2
  CLASS core ;
  FOREIGN XNOR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.9 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.205 0.6 0.695 0.6 0.695 0.53 0.76 0.53 0.76 0.665 0.27 0.665 0.27 0.735 0.205 0.735  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.31 1.315 0.31 1.125 0.375 1.125 0.375 1.315 1.41 1.315 1.41 1.125 1.475 1.125 1.475 1.315 1.9 1.315 1.9 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.9 -0.085 1.9 0.085 1.575 0.085 1.575 0.15 1.51 0.15 1.51 0.365 1.445 0.365 1.445 0.085 0.3 0.085 0.3 0.36 0.235 0.36 0.235 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.355 0.4 0.49 0.4 0.49 0.535 0.355 0.535  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.595 0.335 1.695 0.335 1.695 1.065 1.595 1.065  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.555 0.86 0.62 0.86 0.62 1.155 0.555 1.155  ;
        POLYGON 0.05 0.24 0.115 0.24 0.115 0.8 0.335 0.8 0.335 0.73 0.855 0.73 0.855 0.475 0.92 0.475 0.92 0.795 0.78 0.795 0.78 0.995 0.715 0.995 0.715 0.795 0.4 0.795 0.4 0.865 0.19 0.865 0.19 1.155 0.05 1.155  ;
        POLYGON 1.08 1.055 1.115 1.055 1.115 0.345 1.115 0.28 1.25 0.28 1.25 0.345 1.215 0.345 1.215 0.38 1.18 0.38 1.18 1.055 1.215 1.055 1.215 1.12 1.08 1.12  ;
        POLYGON 0.555 0.15 1.38 0.15 1.38 0.54 1.315 0.54 1.315 0.215 0.62 0.215 0.62 0.535 0.555 0.535  ;
        POLYGON 0.98 1.055 1.015 1.055 1.015 1.185 1.28 1.185 1.28 0.995 1.465 0.995 1.465 0.77 1.53 0.77 1.53 1.06 1.345 1.06 1.345 1.25 0.95 1.25 0.95 1.155 0.915 1.155 0.915 0.86 0.985 0.86 0.985 0.41 0.85 0.41 0.85 0.345 0.815 0.345 0.815 0.28 0.95 0.28 0.95 0.345 1.05 0.345 1.05 0.925 0.98 0.925  ;
  END
END XNOR2_X2

MACRO FILL1  #FILLCELL_X1
  CLASS core ;
  #FOREIGN FILLCELL_X1 0.0 0.0 ;
  FOREIGN FILL1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.19 BY 1.4 ;
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.065 1.315 0.19 1.315 0.19 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.19 -0.085 0.19 0.085 0.065 0.085 0 0.085  ;
    END
  END GRND  #VSS
END FILL1  #FILLCELL_X1

MACRO FILL2  #FILLCELL_X2
  CLASS core ;
  #FOREIGN FILLCELL_X2 0.0 0.0 ;
  FOREIGN FILL2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.065 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0 0.085  ;
    END
  END GRND  #VSS
END FILL2  #FILLCELL_X2

MACRO FILL4  #FILLCELL_X4
  CLASS core ;
  #FOREIGN FILLCELL_X4 0.0 0.0 ;
  FOREIGN FILL4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.065 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0 0.085  ;
    END
  END GRND  #VSS
END FILL4  #FILLCELL_X4

MACRO FILL8  #FILLCELL_X8
  CLASS core ;
  #FOREIGN FILLCELL_X8 0.0 0.0 ;
  FOREIGN FILL8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.065 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 0 0.085  ;
    END
  END GRND  #VSS
END FILL8  #FILLCELL_X8

MACRO FILLCELL_X16
  CLASS core ;
  FOREIGN FILLCELL_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 3.04 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.065 1.315 3.04 1.315 3.04 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 3.04 -0.085 3.04 0.085 0 0.085  ;
    END
  END VSS
END FILLCELL_X16

MACRO FILLCELL_X32
  CLASS core ;
  FOREIGN FILLCELL_X32 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 6.08 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.065 1.315 6.08 1.315 6.08 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 6.08 -0.085 6.08 0.085 0 0.085  ;
    END
  END VSS
END FILLCELL_X32

MACRO ANTENNA_X1
  CLASS core ;
  FOREIGN ANTENNA_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.04 0.42 0.175 0.42 0.175 0.76 0.04 0.76  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.065 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0.065 0.085 0 0.085  ;
    END
  END VSS
END ANTENNA_X1

MACRO LOGIC0_X1
  CLASS core ;
  FOREIGN LOGIC0_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.07 0.265 0.17 0.265 0.17 0.4 0.07 0.4  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.105 1.315 0.105 0.81 0.17 0.81 0.17 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0.17 0.085 0.17 0.2 0.135 0.2 0.07 0.2 0.07 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER M1 ;
        POLYGON 0.085 0.66 0.12 0.66 0.12 0.465 0.22 0.465 0.22 0.725 0.085 0.725  ;
  END
END LOGIC0_X1

MACRO LOGIC1_X1
  CLASS core ;
  FOREIGN LOGIC1_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.07 0.825 0.17 0.825 0.17 0.96 0.07 0.96  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.105 1.315 0.105 1.025 0.17 1.025 0.17 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0.215 0.085 0.215 0.37 0.15 0.37 0.15 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER M1 ;
        POLYGON 0.13 0.455 0.265 0.455 0.265 0.715 0.165 0.715 0.165 0.555 0.13 0.555  ;
  END
END LOGIC1_X1

MACRO MX2X1  #MUX2_X1
  CLASS core ;
  #FOREIGN MUX2_X1 0.0 0.0 ;
  FOREIGN MX2X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN Y  #Z
    DIRECTION OUTPUT ;
	CAPACITANCE 0.000629 ;
	RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 1.35 0.905 1.42 0.905 1.42 0.54 1.375 0.54 1.375 0.44 1.375 0.38 1.35 0.38 1.35 0.245 1.45 0.245 1.45 0.28 1.485 0.28 1.485 1.005 1.45 1.005 1.45 1.04 1.35 1.04  ;
    END
  END Y  #Z
  PIN S0  #S
    DIRECTION INPUT ;
	CAPACITANCE 0.000928 ;
	RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.215 0.545 0.35 0.545 0.35 0.68 0.215 0.68  ;
    END
  END S0  #S
  PIN B  #A
    DIRECTION INPUT ;
	CAPACITANCE 0.000952 ;
	RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.6 0.445 0.665 0.445 0.665 0.48 0.7 0.48 0.7 0.625 0.805 0.625 0.805 0.58 0.905 0.58 0.905 0.625 1.19 0.625 1.19 0.69 0.635 0.69 0.635 0.58 0.6 0.58  ;
    END
  END B  #A
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.285 1.315 0.285 1.01 0.35 1.01 0.35 1.315 1.17 1.315 1.17 1.01 1.235 1.01 1.235 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 1.265 0.085 1.265 0.15 1.2 0.15 1.2 0.275 1.135 0.275 1.135 0.085 0.365 0.085 0.365 0.275 0.3 0.275 0.3 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN A  #B
    DIRECTION INPUT ;
	CAPACITANCE 0.000629 ;
	RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.995 0.425 1.095 0.425 1.095 0.56 0.995 0.56  ;
    END
  END A  #B
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.245 0.15 0.245 0.15 0.78 0.34 0.78 0.34 0.745 0.405 0.745 0.405 0.88 0.34 0.88 0.34 0.845 0.2 0.845 0.2 1.04 0.05 1.04  ;
        POLYGON 0.495 1.01 0.56 1.01 0.56 1.105 0.985 1.105 0.985 1.01 1.05 1.01 1.05 1.17 0.495 1.17  ;
        POLYGON 0.535 0.81 0.705 0.81 0.705 0.815 1.225 0.815 1.225 0.745 1.29 0.745 1.29 0.88 0.745 0.88 0.745 1.04 0.68 1.04 0.68 0.875 0.47 0.875 0.47 0.28 0.68 0.28 0.68 0.245 0.745 0.245 0.745 0.38 0.68 0.38 0.68 0.345 0.535 0.345  ;
  END
END MX2X1  #MUX2_X1

MACRO MUX2_X2
  CLASS core ;
  FOREIGN MUX2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.35 0.87 1.42 0.87 1.42 0.54 1.375 0.54 1.375 0.44 1.375 0.385 1.35 0.385 1.35 0.25 1.45 0.25 1.45 0.285 1.485 0.285 1.485 1.005 1.45 1.005 1.45 1.145 1.35 1.145  ;
    END
  END Z
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.22 0.545 0.32 0.545 0.32 0.68 0.22 0.68  ;
    END
  END S
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.6 0.445 0.665 0.445 0.665 0.48 0.81 0.48 0.81 0.61 1.09 0.61 1.09 0.575 1.155 0.575 1.155 0.71 1.09 0.71 1.09 0.675 0.745 0.675 0.745 0.545 0.665 0.545 0.665 0.58 0.6 0.58  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.26 1.315 0.26 0.975 0.325 0.975 0.325 1.315 1.2 1.315 1.2 0.925 1.265 0.925 1.265 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 1.165 0.085 1.165 0.15 1.1 0.15 1.1 0.28 1.035 0.28 1.035 0.085 0.34 0.085 0.34 0.28 0.275 0.28 0.275 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.92 0.41 1.02 0.41 1.02 0.545 0.92 0.545  ;
    END
  END B
  OBS
      LAYER M1 ;
        POLYGON 0.04 0.25 0.155 0.25 0.155 0.745 0.415 0.745 0.415 0.81 0.175 0.81 0.175 1.005 0.04 1.005  ;
        POLYGON 0.47 0.975 0.535 0.975 0.535 1.07 0.985 1.07 0.985 0.975 1.05 0.975 1.05 1.135 0.47 1.135  ;
        POLYGON 0.535 0.645 0.68 0.645 0.68 0.78 1.225 0.78 1.225 0.71 1.29 0.71 1.29 0.845 0.72 0.845 0.72 1.005 0.655 1.005 0.655 0.84 0.615 0.84 0.615 0.71 0.47 0.71 0.47 0.28 0.655 0.28 0.655 0.245 0.72 0.245 0.72 0.38 0.655 0.38 0.655 0.345 0.535 0.345  ;
  END
END MUX2_X2

MACRO OAI221_X1
  CLASS core ;
  FOREIGN OAI221_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.545 0.63 0.545 0.63 0.68 0.53 0.68  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.425 1.315 0.425 1.155 0.49 1.155 0.49 1.315 1.01 1.315 1.01 1.155 1.075 1.155 1.075 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.705 0.825 0.805 0.825 0.805 0.96 0.705 0.96  ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.3 1.025 0.695 1.025 0.695 1.165 0.63 1.165 0.63 1.09 0.115 1.09 0.115 1.165 0.05 1.165 0.05 1.025 0.235 1.025 0.235 0.82 0.235 0.72 0.235 0.28 0.3 0.28 0.3 0.72 0.335 0.72 0.335 0.82 0.3 0.82  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.07 0.72 0.17 0.72 0.17 0.855 0.07 0.855  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.885 0.085 0.885 0.32 0.82 0.32 0.82 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.895 0.72 0.995 0.72 0.995 0.855 0.895 0.855  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.44 0.465 0.44 0.465 0.575 0.365 0.575  ;
    END
  END C2
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.15 0.49 0.15 0.49 0.32 0.425 0.32 0.425 0.215 0.115 0.215 0.115 0.32 0.05 0.32  ;
        POLYGON 0.635 0.28 0.7 0.28 0.7 0.385 1.01 0.385 1.01 0.28 1.075 0.28 1.075 0.45 0.635 0.45  ;
  END
END OAI221_X1

MACRO OAI221_X2
  CLASS core ;
  FOREIGN OAI221_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.58 0.63 0.58 0.63 0.715 0.53 0.715  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.425 1.315 0.425 1.025 0.49 1.025 0.49 1.315 1.01 1.315 1.01 1.025 1.075 1.025 1.075 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.705 0.685 0.805 0.685 0.805 0.82 0.705 0.82  ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.3 0.885 0.695 0.885 0.695 1.16 0.63 1.16 0.63 0.95 0.115 0.95 0.115 1.16 0.05 1.16 0.05 0.885 0.235 0.885 0.235 0.54 0.235 0.44 0.235 0.375 0.3 0.375 0.3 0.44 0.335 0.44 0.335 0.54 0.3 0.54  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.07 0.58 0.17 0.58 0.17 0.715 0.07 0.715  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.885 0.085 0.885 0.385 0.82 0.385 0.82 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.895 0.58 0.995 0.58 0.995 0.715 0.895 0.715  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.685 0.465 0.685 0.465 0.82 0.365 0.82  ;
    END
  END C2
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.15 0.49 0.15 0.49 0.285 0.425 0.285 0.425 0.215 0.115 0.215 0.115 0.285 0.05 0.285  ;
        POLYGON 0.635 0.375 0.7 0.375 0.7 0.45 1.01 0.45 1.01 0.375 1.075 0.375 1.075 0.515 0.635 0.515  ;
  END
END OAI221_X2

MACRO OAI221_X4
  CLASS core ;
  FOREIGN OAI221_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.71 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.45 0.685 0.55 0.685 0.55 0.82 0.45 0.82  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.425 1.315 0.425 1.11 0.49 1.11 0.49 1.315 1.02 1.315 1.02 1.11 1.085 1.11 1.085 1.315 1.395 1.315 1.395 1.01 1.46 1.01 1.46 1.315 1.71 1.315 1.71 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.745 0.69 0.845 0.69 0.845 0.825 0.745 0.825  ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.545 0.365 1.58 0.365 1.58 0.225 1.645 0.225 1.645 0.58 1.665 0.58 1.665 0.68 1.645 0.68 1.645 0.96 1.58 0.96 1.58 0.82 1.545 0.82  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.07 0.58 0.17 0.58 0.17 0.715 0.07 0.715  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.71 -0.085 1.71 0.085 1.46 0.085 1.46 0.355 1.395 0.355 1.395 0.085 0.895 0.085 0.895 0.32 0.83 0.32 0.83 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.915 0.825 1.015 0.825 1.015 0.96 0.915 0.96  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.44 0.5 0.44 0.5 0.575 0.365 0.575  ;
    END
  END C2
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.15 0.49 0.15 0.49 0.32 0.425 0.32 0.425 0.215 0.115 0.215 0.115 0.32 0.05 0.32  ;
        POLYGON 0.645 0.28 0.71 0.28 0.71 0.385 1.02 0.385 1.02 0.28 1.085 0.28 1.085 0.45 0.645 0.45  ;
        POLYGON 0.05 0.975 0.235 0.975 0.235 0.28 0.3 0.28 0.3 0.975 0.615 0.975 0.615 0.56 1.08 0.56 1.08 0.525 1.145 0.525 1.145 0.66 1.08 0.66 1.08 0.625 0.68 0.625 0.68 0.985 0.705 0.985 0.705 1.12 0.64 1.12 0.64 1.04 0.115 1.04 0.115 1.12 0.05 1.12  ;
        POLYGON 1.175 0.72 1.21 0.72 1.21 0.465 1.175 0.465 1.175 0.33 1.24 0.33 1.24 0.405 1.275 0.405 1.275 0.56 1.415 0.56 1.415 0.525 1.48 0.525 1.48 0.66 1.415 0.66 1.415 0.625 1.275 0.625 1.275 0.78 1.24 0.78 1.24 0.995 1.175 0.995  ;
  END
END OAI221_X4

MACRO AOI222_X1
  CLASS core ;
  FOREIGN AOI222_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 0.875 0.115 0.875 0.115 1.315 0.425 1.315 0.425 0.875 0.49 0.875 0.49 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.805 0.44 0.905 0.44 0.905 0.575 0.805 0.575  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.98 0.58 1.08 0.58 1.08 0.715 0.98 0.715  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.275 0.44 1.375 0.44 1.375 0.575 1.275 0.575  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.115 0.165 0.18 0.165 0.18 0.31 0.875 0.31 0.875 0.165 0.94 0.165 0.94 0.31 1.21 0.31 1.21 0.72 1.285 0.72 1.285 0.82 1.21 0.82 1.21 1.105 1.145 1.105 1.145 0.375 0.115 0.375  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.15 0.545 0.25 0.545 0.25 0.68 0.15 0.68  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 1.38 0.085 1.38 0.15 1.315 0.15 1.315 0.245 1.25 0.245 1.25 0.085 0.555 0.085 0.555 0.245 0.49 0.245 0.49 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.615 0.545 0.715 0.545 0.715 0.68 0.615 0.68  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.35 0.44 0.45 0.44 0.45 0.575 0.35 0.575  ;
    END
  END C2
  OBS
      LAYER M1 ;
        POLYGON 0.24 0.745 0.83 0.745 0.83 1.105 0.765 1.105 0.765 0.81 0.305 0.81 0.305 1.105 0.24 1.105  ;
        POLYGON 0.58 0.875 0.645 0.875 0.645 1.17 0.955 1.17 0.955 0.875 1.02 0.875 1.02 1.17 1.335 1.17 1.335 0.875 1.4 0.875 1.4 1.235 0.58 1.235  ;
  END
END AOI222_X1

MACRO AOI222_X2
  CLASS core ;
  FOREIGN AOI222_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.045 0.115 1.045 0.115 1.315 0.425 1.315 0.425 1.045 0.49 1.045 0.49 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.805 0.58 0.905 0.58 0.905 0.715 0.805 0.715  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.98 0.58 1.08 0.58 1.08 0.715 0.98 0.715  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.275 0.545 1.375 0.545 1.375 0.68 1.275 0.68  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.115 0.155 0.18 0.155 0.18 0.45 0.875 0.45 0.875 0.155 0.94 0.155 0.94 0.45 1.21 0.45 1.21 1.015 1.145 1.015 1.145 0.515 0.115 0.515  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.15 0.58 0.25 0.58 0.25 0.715 0.15 0.715  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 1.38 0.085 1.38 0.15 1.315 0.15 1.315 0.385 1.25 0.385 1.25 0.085 0.555 0.085 0.555 0.385 0.49 0.385 0.49 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.615 0.58 0.715 0.58 0.715 0.715 0.615 0.715  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.35 0.58 0.45 0.58 0.45 0.715 0.35 0.715  ;
    END
  END C2
  OBS
      LAYER M1 ;
        POLYGON 0.24 0.78 0.83 0.78 0.83 1.055 0.765 1.055 0.765 0.845 0.305 0.845 0.305 1.055 0.24 1.055  ;
        POLYGON 0.58 0.91 0.645 0.91 0.645 1.12 0.955 1.12 0.955 0.91 1.02 0.91 1.02 1.12 1.335 1.12 1.335 0.91 1.4 0.91 1.4 1.185 0.58 1.185  ;
  END
END AOI222_X2

MACRO AOI222_X4
  CLASS core ;
  FOREIGN AOI222_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 2.09 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 0.875 0.115 0.875 0.115 1.315 0.425 1.315 0.425 0.875 0.49 0.875 0.49 1.315 1.735 1.315 1.735 1 1.8 1 1.8 1.315 2.09 1.315 2.09 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.805 0.44 0.905 0.44 0.905 0.575 0.805 0.575  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.975 0.58 1.11 0.58 1.11 0.715 0.975 0.715  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.305 0.655 1.405 0.655 1.405 0.79 1.305 0.79  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.885 0.355 1.92 0.355 1.92 0.215 1.985 0.215 1.985 0.3 2.045 0.3 2.045 0.4 1.985 0.4 1.985 0.95 1.92 0.95 1.92 0.81 1.885 0.81  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.15 0.545 0.25 0.545 0.25 0.68 0.15 0.68  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 2.09 -0.085 2.09 0.085 1.8 0.085 1.8 0.345 1.735 0.345 1.735 0.085 1.335 0.085 1.335 0.245 1.27 0.245 1.27 0.085 0.555 0.085 0.555 0.245 0.49 0.245 0.49 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.615 0.545 0.715 0.545 0.715 0.68 0.615 0.68  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.35 0.44 0.45 0.44 0.45 0.575 0.35 0.575  ;
    END
  END C2
  OBS
      LAYER M1 ;
        POLYGON 0.24 0.745 0.83 0.745 0.83 1.105 0.765 1.105 0.765 0.81 0.305 0.81 0.305 1.105 0.24 1.105  ;
        POLYGON 0.115 0.165 0.18 0.165 0.18 0.31 0.895 0.31 0.895 0.165 0.96 0.165 0.96 0.31 1.24 0.31 1.24 0.525 1.36 0.525 1.36 0.455 1.425 0.455 1.425 0.59 1.24 0.59 1.24 1.105 1.175 1.105 1.175 0.375 0.115 0.375  ;
        POLYGON 0.58 0.875 0.645 0.875 0.645 1.17 0.955 1.17 0.955 0.875 1.02 0.875 1.02 1.17 1.36 1.17 1.36 0.875 1.425 0.875 1.425 1.235 0.58 1.235  ;
        POLYGON 1.515 0.355 1.58 0.355 1.58 0.55 1.755 0.55 1.755 0.515 1.82 0.515 1.82 0.65 1.755 0.65 1.755 0.615 1.58 0.615 1.58 0.95 1.515 0.95  ;
  END
END AOI222_X4

MACRO AND2X1  #AND2_X1
  CLASS core ;
  #FOREIGN AND2_X1 0.0 0.0 ;
  FOREIGN AND2X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.25 1.315 0.25 0.95 0.315 0.95 0.315 1.315 0.645 1.315 0.645 0.95 0.71 0.95 0.71 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN A  #A1
    DIRECTION INPUT ;
	CAPACITANCE 0.000603 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.48 0.565 0.58 0.565 0.58 0.7 0.48 0.7  ;
    END
  END A  #A1
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.335 0.085 0.335 0.36 0.27 0.36 0.27 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN B  #A2
    DIRECTION INPUT ;
	CAPACITANCE 0.000411 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.285 0.44 0.42 0.44 0.42 0.54 0.285 0.54  ;
    END
  END B  #A2
  PIN Y  #ZN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
	RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.89 0.085 0.89 0.085 0.54 0.045 0.54 0.045 0.44 0.05 0.44 0.05 0.415 0.05 0.28 0.115 0.28 0.115 0.315 0.15 0.315 0.15 0.99 0.115 0.99 0.115 1.025 0.05 1.025  ;
    END
  END Y #ZN
  OBS
      LAYER M1 ;
        POLYGON 0.215 0.73 0.28 0.73 0.28 0.765 0.645 0.765 0.645 0.28 0.71 0.28 0.71 0.83 0.525 0.83 0.525 1.025 0.46 1.025 0.46 0.83 0.28 0.83 0.28 0.865 0.215 0.865  ;
  END
END AND2X1  #AND2_X1

MACRO AND2_X2
  CLASS core ;
  FOREIGN AND2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 0.925 0.3 0.925 0.3 1.315 0.645 1.315 0.645 0.93 0.71 0.93 0.71 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.48 0.545 0.58 0.545 0.58 0.68 0.48 0.68  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.3 0.085 0.3 0.31 0.235 0.31 0.235 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.315 0.44 0.415 0.44 0.415 0.575 0.315 0.575  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.87 0.085 0.87 0.085 0.54 0.045 0.54 0.045 0.44 0.05 0.44 0.05 0.415 0.05 0.28 0.115 0.28 0.115 0.315 0.15 0.315 0.15 1.005 0.115 1.005 0.115 1.145 0.05 1.145  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.215 0.71 0.28 0.71 0.28 0.745 0.645 0.745 0.645 0.28 0.71 0.28 0.71 0.81 0.525 0.81 0.525 1.005 0.46 1.005 0.46 0.81 0.28 0.81 0.28 0.845 0.215 0.845  ;
  END
END AND2_X2

MACRO AND2_X4
  CLASS core ;
  FOREIGN AND2_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 1.06 0.3 1.06 0.3 1.315 0.645 1.315 0.645 1.015 0.71 1.015 0.71 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.48 0.685 0.58 0.685 0.58 0.82 0.48 0.82  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.3 0.085 0.3 0.265 0.235 0.265 0.235 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.34 0.44 0.475 0.44 0.475 0.54 0.34 0.54  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.045 0.58 0.05 0.58 0.05 0.55 0.05 0.275 0.115 0.275 0.115 0.415 0.15 0.415 0.15 0.87 0.115 0.87 0.115 1.01 0.05 1.01 0.05 0.735 0.05 0.68 0.045 0.68  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.215 0.575 0.28 0.575 0.28 0.885 0.645 0.885 0.645 0.185 0.71 0.185 0.71 0.95 0.525 0.95 0.525 1.09 0.46 1.09 0.46 0.95 0.215 0.95  ;
  END
END AND2_X4

MACRO XOR2X1  #XOR2_X1
  CLASS core ;
  #FOREIGN XOR2_X1 0.0 0.0 ;
  FOREIGN XOR2X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN Y  #Z
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
	RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.775 0.88 0.845 0.88 0.845 0.505 0.6 0.505 0.6 0.44 0.91 0.44 0.91 0.945 0.775 0.945  ;
    END
  END Y  #Z
  PIN A
    DIRECTION INPUT ;
	CAPACITANCE 0.001023 ;
	RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.285 0.685 0.385 0.685 0.385 0.82 0.285 0.82  ;
    END
  END A
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.425 1.315 0.425 0.97 0.49 0.97 0.49 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 1.14 0.085 1.14 0.15 1.075 0.15 1.075 0.49 1.01 0.49 1.01 0.085 0.49 0.085 0.49 0.49 0.425 0.49 0.425 0.085 0.115 0.085 0.115 0.49 0.05 0.49 0.05 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN B
    DIRECTION INPUT ;
	CAPACITANCE 0.000922 ;
	RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.68 0.57 0.78 0.57 0.78 0.705 0.68 0.705  ;
    END
  END B
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.555 0.24 0.555 0.24 0.37 0.305 0.37 0.305 0.555 0.555 0.555 0.555 0.69 0.49 0.69 0.49 0.62 0.115 0.62 0.115 0.98 0.05 0.98  ;
        POLYGON 0.62 0.94 0.685 0.94 0.685 1.01 1.01 1.01 1.01 0.94 1.075 0.94 1.075 1.075 0.62 1.075  ;
  END
END XOR2X1  #XOR2_X1

MACRO XOR2_X2
  CLASS core ;
  FOREIGN XOR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.775 0.74 0.81 0.74 0.81 0.705 0.845 0.705 0.845 0.455 0.62 0.455 0.62 0.32 0.685 0.32 0.685 0.39 0.805 0.39 0.805 0.3 0.905 0.3 0.905 0.39 0.91 0.39 0.91 0.74 0.91 0.945 0.775 0.945  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.295 0.545 0.395 0.545 0.395 0.68 0.295 0.68  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.425 1.315 0.425 0.885 0.49 0.885 0.49 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 1.125 0.085 1.125 0.15 1.06 0.15 1.06 0.335 0.995 0.335 0.995 0.085 0.49 0.085 0.49 0.35 0.425 0.35 0.425 0.085 0.115 0.085 0.115 0.35 0.05 0.35 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.65 0.545 0.75 0.545 0.75 0.68 0.65 0.68  ;
    END
  END B
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.415 0.235 0.415 0.235 0.32 0.3 0.32 0.3 0.415 0.555 0.415 0.555 0.615 0.49 0.615 0.49 0.48 0.115 0.48 0.115 0.98 0.05 0.98  ;
        POLYGON 0.62 0.8 0.685 0.8 0.685 1.01 0.995 1.01 0.995 0.8 1.06 0.8 1.06 1.075 0.62 1.075  ;
  END
END XOR2_X2

MACRO NOR2X1  #NOR2_X1
  CLASS core ;
  #FOREIGN NOR2_X1 0.0 0.0 ;
  FOREIGN NOR2X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 0.865 0.115 0.865 0.115 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN A  #A1
    DIRECTION INPUT ;
	CAPACITANCE 0.000742 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.58 0.505 0.58 0.505 0.68 0.37 0.68  ;
    END
  END A  #A1
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.49 0.085 0.49 0.515 0.425 0.515 0.425 0.085 0.115 0.085 0.115 0.515 0.05 0.515 0.05 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN B  #A2
    DIRECTION INPUT ;
	CAPACITANCE 0.000565 ;
	RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.075 0.58 0.175 0.58 0.175 0.715 0.075 0.715  ;
    END
  END B  #A2
  PIN Y  #ZN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
	RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.4 0.305 0.4 0.305 0.745 0.49 0.745 0.49 0.86 0.525 0.86 0.525 0.96 0.425 0.96 0.425 0.88 0.425 0.86 0.425 0.81 0.24 0.81  ;
    END
  END Y  #ZN
END NOR2X1  #NOR2_X1

MACRO NOR2_X2
  CLASS core ;
  FOREIGN NOR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 0.885 0.115 0.885 0.115 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.545 0.47 0.545 0.47 0.68 0.37 0.68  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.49 0.085 0.49 0.31 0.425 0.31 0.425 0.085 0.115 0.085 0.115 0.31 0.05 0.31 0.05 0.15 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.075 0.44 0.175 0.44 0.175 0.575 0.075 0.575  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.28 0.305 0.28 0.305 0.745 0.49 0.745 0.49 0.86 0.525 0.86 0.525 0.96 0.49 0.96 0.49 1.02 0.425 1.02 0.425 0.96 0.425 0.86 0.425 0.81 0.24 0.81  ;
    END
  END ZN
END NOR2_X2

MACRO NOR2_X4
  CLASS core ;
  FOREIGN NOR2_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.615 1.315 0.615 0.885 0.68 0.885 0.68 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.545 0.465 0.545 0.465 0.68 0.365 0.68  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.87 0.085 0.87 0.285 0.805 0.285 0.805 0.085 0.49 0.085 0.49 0.285 0.425 0.285 0.425 0.085 0.115 0.085 0.115 0.285 0.05 0.285 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.74 0.44 0.84 0.44 0.84 0.575 0.74 0.575  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.255 0.3 0.255 0.3 0.35 0.615 0.35 0.615 0.255 0.68 0.255 0.68 0.415 0.3 0.415 0.3 0.98 0.235 0.98  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.835 0.115 0.835 0.115 1.045 0.425 1.045 0.425 0.755 0.87 0.755 0.87 1.03 0.805 1.03 0.805 0.82 0.49 0.82 0.49 1.11 0.05 1.11  ;
  END
END NOR2_X4

MACRO INVX1
  CLASS core ;
  #FOREIGN INV_X1 0.0 0.0 ;
  FOREIGN INVX1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
	CAPACITANCE 0.000637 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.04 0.465 0.14 0.465 0.14 0.6 0.04 0.6  ;
    END
  END A
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.055 1.315 0.055 0.685 0.12 0.685 0.12 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0.115 0.085 0.115 0.16 0.18 0.16 0.18 0.225 0.115 0.225 0.115 0.4 0.05 0.4 0.05 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN Y  #ZN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.205 0.285 0.34 0.285 0.34 0.76 0.205 0.76  ;
    END
  END Y  #ZN
END INVX1  #INV_X1

MACRO INVX2  #INV_X2
  CLASS core ;
  #FOREIGN INV_X2 0.0 0.0 ;
  FOREIGN INVX2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
	CAPACITANCE 0.000415 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.07 0.465 0.17 0.465 0.17 0.6 0.07 0.6  ;
    END
  END A
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 0.68 0.115 0.68 0.115 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0.18 0.085 0.18 0.15 0.115 0.15 0.115 0.335 0.05 0.335 0.05 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN Y  #ZN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.016000 ;
    RESISTANCE 120.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.305 0.335 0.305 0.335 0.9 0.235 0.9  ;
    END
  END Y  #ZN
END INVX2  #INV_X2

MACRO INVX4  #INV_X4
  CLASS core ;
  #FOREIGN INV_X4 0.0 0.0 ;
  FOREIGN INVX4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
	CAPACITANCE 0.000405 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.07 0.545 0.17 0.545 0.17 0.68 0.07 0.68  ;
    END
  END A
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.03 0.115 1.03 0.115 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0.18 0.085 0.18 0.15 0.115 0.15 0.115 0.375 0.05 0.375 0.05 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN Y  #ZN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.032000 ;
    RESISTANCE 60.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.245 0.335 0.245 0.335 0.98 0.235 0.98  ;
    END
  END Y  #ZN
END INVX4  #INV_X4

MACRO INVX8  #INV_X8
  CLASS core ;
  #FOREIGN INV_X8 0.0 0.0 ;
  FOREIGN INVX8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
	CAPACITANCE 0.000702 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.545 0.465 0.545 0.465 0.68 0.365 0.68  ;
    END
  END A
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.03 0.115 1.03 0.115 1.315 0.425 1.315 0.425 1.03 0.49 1.03 0.49 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.49 0.085 0.49 0.375 0.425 0.375 0.425 0.085 0.115 0.085 0.115 0.375 0.05 0.375 0.05 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN Y  #ZN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.064000 ;
    RESISTANCE 30.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.2 0.245 0.3 0.245 0.3 0.98 0.2 0.98  ;
    END
  END Y  #ZN
END INVX8  #INV_X8

MACRO INV_X16
  CLASS core ;
  FOREIGN INV_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.425 0.545 0.525 0.545 0.525 0.68 0.425 0.68  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.03 0.115 1.03 0.115 1.315 0.425 1.315 0.425 1.03 0.49 1.03 0.49 1.315 0.805 1.315 0.805 1.03 0.87 1.03 0.87 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.87 0.085 0.87 0.35 0.805 0.35 0.805 0.085 0.49 0.085 0.49 0.35 0.425 0.35 0.425 0.085 0.115 0.085 0.115 0.35 0.05 0.35 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.205 0.305 0.205 0.305 0.415 0.615 0.415 0.615 0.4 0.615 0.3 0.615 0.205 0.68 0.205 0.68 0.3 0.715 0.3 0.715 0.4 0.68 0.4 0.68 0.48 0.305 0.48 0.305 0.745 0.68 0.745 0.68 1.02 0.615 1.02 0.615 0.81 0.305 0.81 0.305 1.02 0.24 1.02  ;
    END
  END ZN
END INV_X16

MACRO INV_X32
  CLASS core ;
  FOREIGN INV_X32 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.71 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.04 0.3 0.175 0.3 0.175 0.435 0.04 0.435  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.425 1.315 0.425 1.03 0.49 1.03 0.49 1.315 0.805 1.315 0.805 1.03 0.87 1.03 0.87 1.315 1.185 1.315 1.185 1.03 1.25 1.03 1.25 1.315 1.565 1.315 1.565 1.03 1.63 1.03 1.63 1.315 1.71 1.315 1.71 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.71 -0.085 1.71 0.085 1.63 0.085 1.63 0.345 1.565 0.345 1.565 0.085 1.25 0.085 1.25 0.345 1.185 0.345 1.185 0.085 0.87 0.085 0.87 0.345 0.805 0.345 0.805 0.085 0.49 0.085 0.49 0.345 0.425 0.345 0.425 0.085 0 0.085  ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.265 0.305 0.265 0.305 0.63 0.425 0.63 0.425 0.58 0.525 0.58 0.525 0.63 0.615 0.63 0.615 0.265 0.68 0.265 0.68 0.475 0.995 0.475 0.995 0.265 1.06 0.265 1.06 0.475 1.375 0.475 1.375 0.265 1.44 0.265 1.44 0.905 1.375 0.905 1.375 0.54 1.06 0.54 1.06 0.905 0.995 0.905 0.995 0.54 0.68 0.54 0.68 0.905 0.615 0.905 0.615 0.695 0.305 0.695 0.305 0.905 0.24 0.905  ;
    END
  END ZN
END INV_X32

MACRO AOI22X1  #AOI22_X1
  CLASS core ;
  #FOREIGN AOI22_X1 0.0 0.0 ;
  FOREIGN AOI22X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.615 1.315 0.615 1.015 0.68 1.015 0.68 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END POWR #VDD
  PIN B0  #B1
    DIRECTION INPUT ;
	CAPACITANCE 0.000355 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.525 0.44 0.625 0.44 0.625 0.575 0.525 0.575  ;
    END
  END B0  #B1
  PIN A0  #A1
    DIRECTION INPUT ;
	CAPACITANCE 0.000382 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.685 0.47 0.685 0.47 0.82 0.37 0.82  ;
    END
  END A0  #A1
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.87 0.085 0.87 0.36 0.805 0.36 0.805 0.085 0.115 0.085 0.115 0.36 0.05 0.36 0.05 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN B1  #B2
    DIRECTION INPUT ;
	CAPACITANCE 0.000365 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.69 0.545 0.79 0.545 0.79 0.68 0.69 0.68  ;
    END
  END B1  #B2
  PIN A1  #A2
    DIRECTION INPUT ;
	CAPACITANCE 0.000362 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.075 0.58 0.175 0.58 0.175 0.715 0.075 0.715  ;
    END
  END A1  #A2
  PIN Y  #ZN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.3 0.335 0.3 0.335 0.32 0.425 0.32 0.425 0.25 0.49 0.25 0.49 0.385 0.335 0.385 0.335 0.4 0.305 0.4 0.305 1.025 0.24 1.025 0.24 0.4 0.235 0.4  ;
    END
  END Y  #ZN
  OBS
      LAYER M1 ;
        POLYGON 0.05 1.015 0.115 1.015 0.115 1.09 0.43 1.09 0.43 0.885 0.87 0.885 0.87 1.025 0.805 1.025 0.805 0.95 0.495 0.95 0.495 1.155 0.05 1.155  ;
  END
END AOI22X1  #AOI22_X1

MACRO AOI22_X2
  CLASS core ;
  FOREIGN AOI22_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.615 1.315 0.615 0.885 0.68 0.885 0.68 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.535 0.545 0.635 0.545 0.635 0.68 0.535 0.68  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.545 0.47 0.545 0.47 0.68 0.37 0.68  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.87 0.085 0.87 0.475 0.805 0.475 0.805 0.085 0.115 0.085 0.115 0.475 0.05 0.475 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 0.545 0.8 0.545 0.8 0.68 0.7 0.68  ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.075 0.545 0.175 0.545 0.175 0.68 0.075 0.68  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.415 0.425 0.415 0.425 0.4 0.425 0.3 0.425 0.205 0.49 0.205 0.49 0.3 0.525 0.3 0.525 0.4 0.49 0.4 0.49 0.48 0.305 0.48 0.305 0.98 0.24 0.98  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.835 0.115 0.835 0.115 1.045 0.425 1.045 0.425 0.755 0.87 0.755 0.87 1.03 0.805 1.03 0.805 0.82 0.49 0.82 0.49 1.11 0.05 1.11  ;
  END
END AOI22_X2

MACRO AOI22_X4
  CLASS core ;
  FOREIGN AOI22_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.615 1.315 0.615 1.015 0.68 1.015 0.68 1.315 1.21 1.315 1.21 1 1.275 1 1.275 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.535 0.545 0.635 0.545 0.635 0.68 0.535 0.68  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.44 0.47 0.44 0.47 0.575 0.37 0.575  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 1.275 0.085 1.275 0.345 1.21 0.345 1.21 0.085 0.87 0.085 0.87 0.245 0.805 0.245 0.805 0.085 0.115 0.085 0.115 0.245 0.05 0.245 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.7 0.685 0.8 0.685 0.8 0.82 0.7 0.82  ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.075 0.72 0.175 0.72 0.175 0.855 0.075 0.855  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.36 0.355 1.395 0.355 1.395 0.215 1.46 0.215 1.46 0.95 1.395 0.95 1.395 0.81 1.36 0.81  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.05 1.015 0.115 1.015 0.115 1.09 0.43 1.09 0.43 0.885 0.87 0.885 0.87 1.025 0.805 1.025 0.805 0.95 0.495 0.95 0.495 1.155 0.05 1.155  ;
        POLYGON 0.24 0.31 0.43 0.31 0.43 0.165 0.495 0.165 0.495 0.31 0.925 0.31 0.925 0.63 0.86 0.63 0.86 0.375 0.305 0.375 0.305 1.025 0.24 1.025  ;
        POLYGON 0.99 0.675 1.025 0.675 1.025 0.49 0.99 0.49 0.99 0.355 1.055 0.355 1.055 0.39 1.09 0.39 1.09 0.55 1.23 0.55 1.23 0.515 1.295 0.515 1.295 0.65 1.23 0.65 1.23 0.615 1.09 0.615 1.09 0.81 1.055 0.81 1.055 0.95 0.99 0.95  ;
  END
END AOI22_X4

MACRO OAI22X1  #OAI22_X1
  CLASS core ;
  #FOREIGN OAI22_X1 0.0 0.0 ;
  FOREIGN OAI22X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.11 0.115 1.11 0.115 1.315 0.805 1.315 0.805 1.11 0.87 1.11 0.87 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN B0  #B1
    DIRECTION INPUT ;
	CAPACITANCE 0.000356 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.685 0.63 0.685 0.63 0.82 0.53 0.82  ;
    END
  END B0  #B1
  PIN A0  #A1
    DIRECTION INPUT ;
	CAPACITANCE 0.000420 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.555 0.465 0.555 0.465 0.69 0.365 0.69  ;
    END
  END A0  #A1
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.68 0.085 0.68 0.36 0.615 0.36 0.615 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN B1  #B2
    DIRECTION INPUT ;
	CAPACITANCE 0.000357 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.695 0.825 0.795 0.825 0.795 0.96 0.695 0.96  ;
    END
  END B1  #B2
  PIN A1  #A2
    DIRECTION INPUT ;
	CAPACITANCE 0.000420 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.07 0.44 0.17 0.44 0.17 0.575 0.07 0.575  ;
    END
  END A1  #A2
  PIN Y  #ZN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.28 0.3 0.28 0.3 0.875 0.49 0.875 0.49 1.12 0.425 1.12 0.425 0.94 0.235 0.94  ;
    END
  END Y  #ZN
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.15 0.49 0.15 0.49 0.425 0.805 0.425 0.805 0.28 0.87 0.28 0.87 0.49 0.425 0.49 0.425 0.215 0.115 0.215 0.115 0.36 0.05 0.36  ;
  END
END OAI22X1  #OAI22_X1

MACRO OAI22_X2
  CLASS core ;
  FOREIGN OAI22_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.045 0.115 1.045 0.115 1.315 0.805 1.315 0.805 1.045 0.87 1.045 0.87 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.705 0.63 0.705 0.63 0.84 0.53 0.84  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.705 0.465 0.705 0.465 0.84 0.365 0.84  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.68 0.085 0.68 0.51 0.615 0.51 0.615 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.695 0.705 0.795 0.705 0.795 0.84 0.695 0.84  ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.07 0.58 0.17 0.58 0.17 0.715 0.07 0.715  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.28 0.3 0.28 0.3 0.905 0.49 0.905 0.49 1 0.525 1 0.525 1.1 0.49 1.1 0.49 1.18 0.425 1.18 0.425 1.1 0.425 1 0.425 0.97 0.235 0.97  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.15 0.49 0.15 0.49 0.575 0.805 0.575 0.805 0.28 0.87 0.28 0.87 0.64 0.425 0.64 0.425 0.215 0.115 0.215 0.115 0.51 0.05 0.51  ;
  END
END OAI22_X2

MACRO OAI22_X4
  CLASS core ;
  FOREIGN OAI22_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.2 0.115 1.2 0.115 1.315 0.83 1.315 0.83 1.2 0.895 1.2 0.895 1.315 1.19 1.315 1.19 1.04 1.255 1.04 1.255 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.555 0.915 0.69 0.915 0.69 1.05 0.555 1.05  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.26 0.725 0.36 0.725 0.36 0.86 0.26 0.86  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 1.255 0.085 1.255 0.385 1.19 0.385 1.19 0.085 0.705 0.085 0.705 0.4 0.64 0.4 0.64 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.725 0.725 0.825 0.725 0.825 0.86 0.725 0.86  ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.075 0.48 0.175 0.48 0.175 0.615 0.075 0.615  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.375 0.255 1.475 0.255 1.475 0.99 1.375 0.99  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.19 0.52 0.19 0.52 0.465 0.83 0.465 0.83 0.32 0.895 0.32 0.895 0.53 0.455 0.53 0.455 0.255 0.115 0.255 0.115 0.4 0.05 0.4  ;
        POLYGON 0.24 0.32 0.305 0.32 0.305 0.595 0.985 0.595 0.985 0.66 0.49 0.66 0.49 1.21 0.425 1.21 0.425 0.66 0.24 0.66  ;
        POLYGON 0.985 0.725 1.05 0.725 1.05 0.53 0.985 0.53 0.985 0.395 1.05 0.395 1.05 0.43 1.115 0.43 1.115 0.59 1.245 0.59 1.245 0.555 1.31 0.555 1.31 0.69 1.245 0.69 1.245 0.655 1.115 0.655 1.115 0.86 1.05 0.86 1.05 1 0.985 1  ;
  END
END OAI22_X4

MACRO NAND4X1  #NAND4_X1
  CLASS core ;
  #FOREIGN NAND4_X1 0.0 0.0 ;
  FOREIGN NAND4X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.155 0.115 1.155 0.115 1.315 0.425 1.315 0.425 1.155 0.49 1.155 0.49 1.315 0.805 1.315 0.805 1.155 0.87 1.155 0.87 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN C  #A3
    DIRECTION INPUT ;
	CAPACITANCE 0.000368 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.44 0.6 0.44 0.6 0.575 0.5 0.575  ;
    END
  END C  #A3
  PIN A  #A1
    DIRECTION INPUT ;
	CAPACITANCE 0.000403 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.18 0.685 0.28 0.685 0.28 0.82 0.18 0.82  ;
    END
  END A  #A1
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.87 0.085 0.87 0.275 0.805 0.275 0.805 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN B  #A2
    DIRECTION INPUT ;
	CAPACITANCE 0.000545 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.345 0.825 0.445 0.825 0.445 0.96 0.345 0.96  ;
    END
  END B  #A2
  PIN D  #A4
    DIRECTION INPUT ;
	CAPACITANCE 0.000371 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.58 0.8 0.58 0.8 0.715 0.665 0.715  ;
    END
  END D  #A4
  PIN Y  #ZN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.28 0.115 0.28 0.115 1.025 0.615 1.025 0.615 1 0.715 1 0.715 1.1 0.68 1.1 0.68 1.23 0.615 1.23 0.615 1.1 0.615 1.09 0.305 1.09 0.305 1.23 0.24 1.23 0.24 1.09 0.05 1.09  ;
    END
  END Y  #ZN
END NAND4X1  #NAND4_X1

MACRO NAND4_X2
  CLASS core ;
  FOREIGN NAND4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.015 0.115 1.015 0.115 1.315 0.425 1.315 0.425 1.015 0.49 1.015 0.49 1.315 0.815 1.315 0.815 1.015 0.88 1.015 0.88 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.51 0.58 0.61 0.58 0.61 0.715 0.51 0.715  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.18 0.58 0.28 0.58 0.28 0.715 0.18 0.715  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.88 0.085 0.88 0.345 0.815 0.345 0.815 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.345 0.685 0.445 0.685 0.445 0.82 0.345 0.82  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.675 0.685 0.81 0.685 0.81 0.82 0.675 0.82  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.28 0.115 0.28 0.115 0.885 0.68 0.885 0.68 1.235 0.615 1.235 0.615 0.95 0.335 0.95 0.335 1 0.335 1.1 0.3 1.1 0.3 1.235 0.235 1.235 0.235 1.1 0.235 1 0.235 0.95 0.05 0.95  ;
    END
  END ZN
END NAND4_X2

MACRO NAND4_X4
  CLASS core ;
  FOREIGN NAND4_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.9 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.08 1.315 0.08 1.06 0.145 1.06 0.145 1.315 0.42 1.315 0.42 1.235 0.555 1.235 0.555 1.315 0.8 1.315 0.8 1.235 0.935 1.235 0.935 1.315 1.18 1.315 1.18 1.235 1.315 1.235 1.315 1.315 1.56 1.315 1.56 1.235 1.695 1.235 1.695 1.315 1.9 1.315 1.9 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.565 0.715 1.175 0.715 1.175 0.85 1.11 0.85 1.11 0.78 0.63 0.78 0.63 0.85 0.565 0.85  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.185 0.455 1.525 0.455 1.525 0.715 1.46 0.715 1.46 0.52 0.25 0.52 0.25 0.715 0.185 0.715  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.9 -0.085 1.9 0.085 1.715 0.085 1.715 0.26 1.58 0.26 1.58 0.085 0.115 0.085 0.115 0.34 0.05 0.34 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.375 0.585 1.365 0.585 1.365 0.72 1.3 0.72 1.3 0.65 0.44 0.65 0.44 0.72 0.375 0.72  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.695 0.845 0.795 0.845 0.795 0.98 0.695 0.98  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.27 1.045 0.425 1.045 0.425 1 0.525 1 0.525 1.045 1.59 1.045 1.59 0.39 1.46 0.39 1.46 0.355 0.94 0.355 0.94 0.39 0.805 0.39 0.805 0.325 0.84 0.325 0.84 0.29 1.52 0.29 1.52 0.325 1.655 0.325 1.655 1.11 1.47 1.11 1.47 1.18 1.405 1.18 1.405 1.11 1.09 1.11 1.09 1.18 1.025 1.18 1.025 1.11 0.71 1.11 0.71 1.18 0.645 1.18 0.645 1.11 0.335 1.11 0.335 1.18 0.27 1.18  ;
    END
  END ZN
END NAND4_X4

MACRO OR3_X1
  CLASS core ;
  FOREIGN OR3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.27 1.315 0.27 1.015 0.335 1.015 0.335 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.345 0.58 0.445 0.58 0.445 0.715 0.345 0.715  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.72 0.58 0.82 0.58 0.82 0.715 0.72 0.715  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.71 0.085 0.71 0.35 0.645 0.35 0.645 0.085 0.315 0.085 0.315 0.35 0.25 0.35 0.25 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.685 0.63 0.685 0.63 0.82 0.53 0.82  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.97 0.085 0.97 0.085 0.54 0.045 0.54 0.045 0.44 0.085 0.44 0.085 0.37 0.05 0.37 0.05 0.235 0.115 0.235 0.115 0.27 0.15 0.27 0.15 1.07 0.115 1.07 0.115 1.105 0.05 1.105  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.28 0.885 0.9 0.885 0.9 1.245 0.835 1.245 0.835 0.95 0.215 0.95 0.215 0.415 0.28 0.415 0.28 0.45 0.46 0.45 0.46 0.235 0.525 0.235 0.525 0.45 0.835 0.45 0.835 0.235 0.9 0.235 0.9 0.515 0.28 0.515  ;
  END
END OR3_X1

MACRO OR3_X2
  CLASS core ;
  FOREIGN OR3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 1.015 0.3 1.015 0.3 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.345 0.58 0.445 0.58 0.445 0.715 0.345 0.715  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.72 0.58 0.82 0.58 0.82 0.715 0.72 0.715  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.71 0.085 0.71 0.37 0.645 0.37 0.645 0.085 0.3 0.085 0.3 0.285 0.235 0.285 0.235 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.685 0.63 0.685 0.63 0.82 0.53 0.82  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.96 0.085 0.96 0.085 0.54 0.045 0.54 0.045 0.44 0.05 0.44 0.05 0.39 0.05 0.255 0.115 0.255 0.115 0.29 0.15 0.29 0.15 1.095 0.115 1.095 0.115 1.235 0.05 1.235  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.28 0.885 0.9 0.885 0.9 1.235 0.835 1.235 0.835 0.95 0.215 0.95 0.215 0.415 0.28 0.415 0.28 0.45 0.46 0.45 0.46 0.255 0.525 0.255 0.525 0.45 0.835 0.45 0.835 0.255 0.9 0.255 0.9 0.515 0.28 0.515  ;
  END
END OR3_X2

MACRO OR3_X4
  CLASS core ;
  FOREIGN OR3_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.2 1.315 0.2 1.18 0.335 1.18 0.335 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.345 0.685 0.445 0.685 0.445 0.82 0.345 0.82  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.72 0.685 0.82 0.685 0.82 0.82 0.72 0.82  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.71 0.085 0.71 0.475 0.645 0.475 0.645 0.085 0.3 0.085 0.3 0.35 0.235 0.35 0.235 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.685 0.63 0.685 0.63 0.82 0.53 0.82  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.045 0.58 0.085 0.58 0.085 0.495 0.05 0.495 0.05 0.22 0.115 0.22 0.115 0.36 0.15 0.36 0.15 0.815 0.115 0.815 0.115 0.955 0.05 0.955 0.05 0.68 0.045 0.68  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.28 0.885 0.9 0.885 0.9 1.16 0.835 1.16 0.835 0.95 0.215 0.95 0.215 0.52 0.28 0.52 0.28 0.555 0.46 0.555 0.46 0.36 0.525 0.36 0.525 0.555 0.835 0.555 0.835 0.36 0.9 0.36 0.9 0.62 0.28 0.62  ;
  END
END OR3_X4

MACRO AOI21X1  #AOI21_X1
  CLASS core ;
  #FOREIGN AOI21_X1 0.0 0.0 ;
  FOREIGN AOI21X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN A0  #A
    DIRECTION INPUT ;
	CAPACITANCE 0.000347 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.58 0.58 0.715 0.58 0.715 0.715 0.58 0.715  ;
    END
  END A0  #A
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.645 1.315 0.645 0.97 0.71 0.97 0.71 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN A1  #B1
    DIRECTION INPUT ;
	CAPACITANCE 0.000392 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.685 0.505 0.685 0.505 0.82 0.37 0.82  ;
    END
  END A1  #B1
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.71 0.085 0.71 0.395 0.645 0.395 0.645 0.085 0.12 0.085 0.12 0.36 0.055 0.36 0.055 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN B0  #B2
    DIRECTION INPUT ;
	CAPACITANCE 0.000410 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.075 0.44 0.175 0.44 0.175 0.575 0.075 0.575  ;
    END
  END B0  #B2
  PIN Y  #ZN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.3 0.335 0.3 0.335 0.35 0.43 0.35 0.43 0.28 0.495 0.28 0.495 0.415 0.305 0.415 0.305 0.98 0.24 0.98 0.24 0.4 0.235 0.4  ;
    END
  END Y  #ZN
  OBS
      LAYER M1 ;
        POLYGON 0.055 0.97 0.12 0.97 0.12 1.045 0.43 1.045 0.43 0.97 0.495 0.97 0.495 1.11 0.055 1.11  ;
  END
END AOI21X1  #AOI21_X1

MACRO AOI21_X2
  CLASS core ;
  FOREIGN AOI21_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.535 0.545 0.635 0.545 0.635 0.68 0.535 0.68  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.615 1.315 0.615 0.885 0.68 0.885 0.68 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.545 0.47 0.545 0.47 0.68 0.37 0.68  ;
    END
  END B1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.695 0.085 0.695 0.415 0.63 0.415 0.63 0.085 0.115 0.085 0.115 0.475 0.05 0.475 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.075 0.545 0.175 0.545 0.175 0.68 0.075 0.68  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.415 0.425 0.415 0.425 0.4 0.425 0.3 0.425 0.205 0.49 0.205 0.49 0.3 0.525 0.3 0.525 0.4 0.49 0.4 0.49 0.48 0.305 0.48 0.305 0.98 0.24 0.98  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.835 0.115 0.835 0.115 1.045 0.425 1.045 0.425 0.835 0.49 0.835 0.49 1.11 0.05 1.11  ;
  END
END AOI21_X2

MACRO AOI21_X4
  CLASS core ;
  FOREIGN AOI21_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.475 0.735 0.575 0.735 0.575 0.87 0.475 0.87  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.615 1.315 0.615 1.02 0.68 1.02 0.68 1.315 0.99 1.315 0.99 1 1.055 1 1.055 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.31 0.405 0.41 0.405 0.41 0.54 0.31 0.54  ;
    END
  END B1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 1.055 0.085 1.055 0.345 0.99 0.345 0.99 0.085 0.68 0.085 0.68 0.325 0.615 0.325 0.615 0.085 0.115 0.085 0.115 0.325 0.05 0.325 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.08 0.44 0.18 0.44 0.18 0.575 0.08 0.575  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.14 0.355 1.175 0.355 1.175 0.215 1.24 0.215 1.24 0.3 1.285 0.3 1.285 0.4 1.24 0.4 1.24 0.95 1.175 0.95 1.175 0.81 1.14 0.81  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.05 1.02 0.115 1.02 0.115 1.095 0.425 1.095 0.425 1.02 0.49 1.02 0.49 1.16 0.05 1.16  ;
        POLYGON 0.24 0.605 0.475 0.605 0.475 0.34 0.43 0.34 0.43 0.205 0.495 0.205 0.495 0.275 0.54 0.275 0.54 0.515 0.74 0.515 0.74 0.65 0.675 0.65 0.675 0.58 0.54 0.58 0.54 0.67 0.305 0.67 0.305 1.03 0.24 1.03  ;
        POLYGON 0.77 0.71 0.805 0.71 0.805 0.455 0.77 0.455 0.77 0.32 0.835 0.32 0.835 0.355 0.87 0.355 0.87 0.55 1.01 0.55 1.01 0.515 1.075 0.515 1.075 0.65 1.01 0.65 1.01 0.615 0.87 0.615 0.87 0.845 0.835 0.845 0.835 0.985 0.77 0.985  ;
  END
END AOI21_X4

MACRO NOR3X1  #NOR3_X1
  CLASS core ;
  #FOREIGN NOR3_X1 0.0 0.0 ;
  FOREIGN NOR3X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.615 1.315 0.615 0.89 0.68 0.89 0.68 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN C  #A3
    DIRECTION INPUT ;
	CAPACITANCE 0.000502 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.51 0.685 0.645 0.685 0.645 0.82 0.51 0.82  ;
    END
  END C  #A3
  PIN A  #A1
    DIRECTION INPUT ;
	CAPACITANCE 0.000400 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.18 0.685 0.28 0.685 0.28 0.82 0.18 0.82  ;
    END
  END A  #A1
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.68 0.085 0.68 0.385 0.615 0.385 0.615 0.085 0.3 0.085 0.3 0.385 0.235 0.385 0.235 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN B  #A2
    DIRECTION INPUT ;
	CAPACITANCE 0.000564 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.345 0.58 0.445 0.58 0.445 0.715 0.345 0.715  ;
    END
  END B  #A2
  PIN Y  #ZN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.27 0.115 0.27 0.115 0.45 0.425 0.45 0.425 0.27 0.49 0.27 0.49 0.515 0.115 0.515 0.115 1.12 0.05 1.12  ;
    END
  END Y  #ZN
END NOR3X1  #NOR3_X1

MACRO NOR3_X2
  CLASS core ;
  FOREIGN NOR3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.615 1.315 0.615 1.01 0.68 1.01 0.68 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.535 0.44 0.635 0.44 0.635 0.575 0.535 0.575  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.18 0.44 0.28 0.44 0.28 0.575 0.18 0.575  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.68 0.085 0.68 0.245 0.615 0.245 0.615 0.085 0.3 0.085 0.3 0.245 0.235 0.245 0.235 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.345 0.545 0.445 0.545 0.445 0.68 0.345 0.68  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.215 0.115 0.215 0.115 0.31 0.425 0.31 0.425 0.215 0.49 0.215 0.49 0.375 0.115 0.375 0.115 0.98 0.05 0.98  ;
    END
  END ZN
END NOR3_X2

MACRO NOR3_X4
  CLASS core ;
  FOREIGN NOR3_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0.14 1.315 1.21 1.315 1.21 0.96 1.275 0.96 1.275 1.315 1.33 1.315 1.33 1.485 0 1.485 0 1.315 0.075 1.315 0.075 1.2 0.04 1.2 0.04 0.995 0.175 0.995 0.175 1.2 0.14 1.2  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.21 0.495 0.275 0.495 0.275 0.735 1.105 0.735 1.105 0.495 1.17 0.495 1.17 0.8 0.21 0.8  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.495 0.435 0.495 0.435 0.605 0.915 0.605 0.915 0.495 0.98 0.495 0.98 0.67 0.37 0.67  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 1.275 0.085 1.275 0.245 1.21 0.245 1.21 0.085 0.93 0.085 0.93 0.21 0.795 0.21 0.795 0.085 0.55 0.085 0.55 0.21 0.415 0.21 0.415 0.085 0.175 0.085 0.175 0.21 0.04 0.21 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.615 0.405 0.715 0.405 0.715 0.54 0.615 0.54  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.045 0.44 0.08 0.44 0.08 0.275 0.26 0.275 0.26 0.205 0.325 0.205 0.325 0.275 0.64 0.275 0.64 0.205 0.705 0.205 0.705 0.275 1.02 0.275 1.02 0.205 1.085 0.205 1.085 0.34 0.145 0.34 0.145 0.44 0.145 0.54 0.145 0.865 0.705 0.865 0.705 0.9 0.74 0.9 0.74 0.965 0.605 0.965 0.605 0.93 0.08 0.93 0.08 0.54 0.045 0.54  ;
    END
  END ZN
END NOR3_X4

MACRO NAND2X1  #NAND2_X1
  CLASS core ;
  #FOREIGN NAND2_X1 0.0 0.0 ;
  FOREIGN NAND2X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1 0.115 1 0.115 1.315 0.425 1.315 0.425 1 0.49 1 0.49 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN A  #A1
    DIRECTION INPUT ;
	CAPACITANCE 0.000451 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.18 0.58 0.28 0.58 0.28 0.715 0.18 0.715  ;
    END
  END A  #A1
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.49 0.085 0.49 0.5 0.425 0.5 0.425 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN B  #A2
    DIRECTION INPUT ;
	CAPACITANCE 0.000339 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.345 0.685 0.445 0.685 0.445 0.82 0.345 0.82  ;
    END
  END B  #A2
  PIN Y  #ZN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.42 0.115 0.42 0.115 0.87 0.3 0.87 0.3 1 0.335 1 0.335 1.1 0.235 1.1 0.235 1.075 0.235 1 0.235 0.935 0.05 0.935  ;
    END
  END Y  #ZN
END NAND2X1  #NAND2_X1

MACRO NAND2X2  #NAND2_X2
  CLASS core ;
  #FOREIGN NAND2_X2 0.0 0.0 ;
  FOREIGN NAND2X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.015 0.115 1.015 0.115 1.315 0.425 1.315 0.425 1.015 0.49 1.015 0.49 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN A  #A1
    DIRECTION INPUT ;
	CAPACITANCE 0.000712 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.18 0.685 0.28 0.685 0.28 0.82 0.18 0.82  ;
    END
  END A  #A1
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.49 0.085 0.49 0.51 0.425 0.51 0.425 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN B  #A2
    DIRECTION INPUT ;
	CAPACITANCE 0.000450 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.345 0.58 0.445 0.58 0.445 0.715 0.345 0.715  ;
    END
  END B  #A2
  PIN Y  #ZN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.016000 ;
    RESISTANCE 120.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.28 0.115 0.28 0.115 0.885 0.3 0.885 0.3 1 0.335 1 0.335 1.1 0.3 1.1 0.3 1.235 0.235 1.235 0.235 1.1 0.235 1 0.235 0.95 0.05 0.95  ;
    END
  END Y  #ZN
END NAND2X2  #NAND2_X2

MACRO NAND2_X4
  CLASS core ;
  FOREIGN NAND2_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 0.92 0.115 0.92 0.115 1.315 0.425 1.315 0.425 0.92 0.49 0.92 0.49 1.315 0.805 1.315 0.805 0.92 0.87 0.92 0.87 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.075 0.58 0.175 0.58 0.175 0.715 0.075 0.715  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.68 0.085 0.68 0.51 0.615 0.51 0.615 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.745 0.705 0.845 0.705 0.845 0.84 0.745 0.84  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.42 0.305 0.42 0.305 0.79 0.68 0.79 0.68 1 0.715 1 0.715 1.1 0.68 1.1 0.68 1.14 0.615 1.14 0.615 1.1 0.615 1 0.615 0.855 0.305 0.855 0.305 1.14 0.24 1.14  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.24 0.49 0.24 0.49 0.575 0.805 0.575 0.805 0.28 0.87 0.28 0.87 0.64 0.425 0.64 0.425 0.305 0.115 0.305 0.115 0.515 0.05 0.515  ;
  END
END NAND2_X4

MACRO OR2X1  #OR2_X1
  CLASS core ;
  #FOREIGN OR2_X1 0.0 0.0 ;
  FOREIGN OR2X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.27 1.315 0.27 1.11 0.335 1.11 0.335 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN A  #A1
    DIRECTION INPUT ;
	CAPACITANCE 0.000896 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.48 0.72 0.58 0.72 0.58 0.855 0.48 0.855  ;
    END
  END A  #A1
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.71 0.085 0.71 0.49 0.645 0.49 0.645 0.085 0.315 0.085 0.315 0.49 0.25 0.49 0.25 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN B  #A2
    DIRECTION INPUT ;
	CAPACITANCE 0.000358 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.315 0.825 0.415 0.825 0.415 0.96 0.315 0.96  ;
    END
  END B  #A2
  PIN Y  #ZN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.985 0.085 0.985 0.085 0.68 0.045 0.68 0.045 0.58 0.085 0.58 0.085 0.51 0.05 0.51 0.05 0.375 0.115 0.375 0.115 0.41 0.15 0.41 0.15 1.085 0.115 1.085 0.115 1.12 0.05 1.12  ;
    END
  END Y  #ZN
  OBS
      LAYER M1 ;
        POLYGON 0.215 0.555 0.28 0.555 0.28 0.59 0.455 0.59 0.455 0.375 0.52 0.375 0.52 0.59 0.71 0.59 0.71 1.12 0.645 1.12 0.645 0.655 0.28 0.655 0.28 0.69 0.215 0.69  ;
  END
END OR2X1  #OR2_X1

MACRO OR2_X2
  CLASS core ;
  FOREIGN OR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 0.9 0.3 0.9 0.3 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.48 0.58 0.58 0.58 0.58 0.715 0.48 0.715  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.71 0.085 0.71 0.37 0.645 0.37 0.645 0.085 0.3 0.085 0.3 0.285 0.235 0.285 0.235 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.315 0.685 0.415 0.685 0.415 0.82 0.315 0.82  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.845 0.085 0.845 0.085 0.54 0.045 0.54 0.045 0.44 0.05 0.44 0.05 0.39 0.05 0.255 0.115 0.255 0.115 0.29 0.15 0.29 0.15 0.98 0.115 0.98 0.115 1.12 0.05 1.12  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.215 0.415 0.28 0.415 0.28 0.45 0.455 0.45 0.455 0.255 0.52 0.255 0.52 0.45 0.71 0.45 0.71 0.98 0.645 0.98 0.645 0.515 0.28 0.515 0.28 0.55 0.215 0.55  ;
  END
END OR2_X2

MACRO OR2_X4
  CLASS core ;
  FOREIGN OR2_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 1.04 0.3 1.04 0.3 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.685 0.63 0.685 0.63 0.82 0.53 0.82  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.71 0.085 0.71 0.475 0.645 0.475 0.645 0.085 0.3 0.085 0.3 0.35 0.235 0.35 0.235 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.345 0.685 0.445 0.685 0.445 0.82 0.345 0.82  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.045 0.58 0.085 0.58 0.085 0.495 0.05 0.495 0.05 0.22 0.115 0.22 0.115 0.36 0.15 0.36 0.15 0.85 0.115 0.85 0.115 0.99 0.05 0.99 0.05 0.715 0.05 0.68 0.045 0.68  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.28 0.91 0.37 0.91 0.37 0.92 0.645 0.92 0.645 0.885 0.71 0.885 0.71 1.02 0.645 1.02 0.645 0.985 0.335 0.985 0.335 0.975 0.215 0.975 0.215 0.52 0.28 0.52 0.28 0.555 0.455 0.555 0.455 0.36 0.52 0.36 0.52 0.62 0.28 0.62  ;
  END
END OR2_X4

MACRO AOI211_X1
  CLASS core ;
  FOREIGN AOI211_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.715 0.545 0.815 0.545 0.815 0.68 0.715 0.68  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.805 1.315 0.805 0.75 0.87 0.75 0.87 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.76 0.085 0.76 0.15 0.695 0.15 0.695 0.35 0.63 0.35 0.63 0.085 0.115 0.085 0.115 0.35 0.05 0.35 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.535 0.545 0.635 0.545 0.635 0.68 0.535 0.68  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.415 0.425 0.415 0.425 0.27 0.49 0.27 0.49 0.415 0.82 0.415 0.82 0.235 0.885 0.235 0.885 0.48 0.305 0.48 0.305 0.98 0.24 0.98  ;
    END
  END ZN
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.075 0.44 0.175 0.44 0.175 0.575 0.075 0.575  ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.545 0.47 0.545 0.47 0.68 0.37 0.68  ;
    END
  END C1
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.75 0.115 0.75 0.115 1.045 0.425 1.045 0.425 0.75 0.49 0.75 0.49 1.11 0.05 1.11  ;
  END
END AOI211_X1

MACRO AOI211_X2
  CLASS core ;
  FOREIGN AOI211_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.715 0.545 0.815 0.545 0.815 0.68 0.715 0.68  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.805 1.315 0.805 1.01 0.87 1.01 0.87 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.695 0.085 0.695 0.215 0.76 0.215 0.76 0.28 0.695 0.28 0.695 0.35 0.63 0.35 0.63 0.085 0.115 0.085 0.115 0.475 0.05 0.475 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.535 0.545 0.635 0.545 0.635 0.68 0.535 0.68  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.415 0.425 0.415 0.425 0.4 0.425 0.3 0.425 0.205 0.49 0.205 0.49 0.3 0.525 0.3 0.525 0.4 0.525 0.415 0.82 0.415 0.82 0.32 0.885 0.32 0.885 0.48 0.305 0.48 0.305 0.98 0.24 0.98  ;
    END
  END ZN
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.075 0.545 0.175 0.545 0.175 0.68 0.075 0.68  ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.545 0.47 0.545 0.47 0.68 0.37 0.68  ;
    END
  END C1
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.835 0.115 0.835 0.115 1.045 0.425 1.045 0.425 0.835 0.49 0.835 0.49 1.11 0.05 1.11  ;
  END
END AOI211_X2

MACRO AOI211_X4
  CLASS core ;
  FOREIGN AOI211_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.705 0.66 0.805 0.66 0.805 0.795 0.705 0.795  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.82 1.315 0.82 0.865 0.885 0.865 0.885 1.315 1.205 1.315 1.205 1 1.27 1 1.27 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 1.27 0.085 1.27 0.345 1.205 0.345 1.205 0.085 0.695 0.085 0.695 0.27 0.63 0.27 0.63 0.085 0.115 0.085 0.115 0.27 0.05 0.27 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.515 0.465 0.615 0.465 0.615 0.6 0.515 0.6  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.355 0.355 1.39 0.355 1.39 0.215 1.455 0.215 1.455 0.95 1.39 0.95 1.39 0.81 1.355 0.81  ;
    END
  END ZN
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.09 0.58 0.19 0.58 0.19 0.715 0.09 0.715  ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.385 0.66 0.485 0.66 0.485 0.795 0.385 0.795  ;
    END
  END C1
  OBS
      LAYER M1 ;
        POLYGON 0.065 0.865 0.13 0.865 0.13 1.16 0.44 1.16 0.44 0.865 0.505 0.865 0.505 1.225 0.065 1.225  ;
        POLYGON 0.255 0.335 0.425 0.335 0.425 0.19 0.49 0.19 0.49 0.335 0.82 0.335 0.82 0.155 0.92 0.155 0.92 0.515 0.955 0.515 0.955 0.65 0.89 0.65 0.89 0.615 0.855 0.615 0.855 0.4 0.32 0.4 0.32 1.095 0.255 1.095  ;
        POLYGON 0.985 0.71 1.02 0.71 1.02 0.455 0.985 0.455 0.985 0.32 1.05 0.32 1.05 0.355 1.085 0.355 1.085 0.55 1.225 0.55 1.225 0.515 1.29 0.515 1.29 0.65 1.225 0.65 1.225 0.615 1.085 0.615 1.085 0.845 1.05 0.845 1.05 0.985 0.985 0.985  ;
  END
END AOI211_X4

MACRO CLKBUFX1
  CLASS core ;
  FOREIGN CLKBUFX1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN Y  #Z
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.845 0.085 0.845 0.085 0.54 0.045 0.54 0.045 0.44 0.05 0.44 0.05 0.305 0.115 0.305 0.115 0.34 0.15 0.34 0.15 0.945 0.115 0.945 0.115 0.98 0.05 0.98  ;
    END
  END Y  #Z
  PIN A
    DIRECTION INPUT ;
	CAPACITANCE 0.000669 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.255 0.685 0.39 0.685 0.39 0.82 0.255 0.82  ;
    END
  END A
  PIN POWR #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 0.905 0.3 0.905 0.3 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.3 0.085 0.3 0.42 0.235 0.42 0.235 0.085 0 0.085  ;
    END
  END GRND  #VSS
  OBS
      LAYER M1 ;
        POLYGON 0.215 0.485 0.28 0.485 0.28 0.52 0.455 0.52 0.455 0.305 0.52 0.305 0.52 0.98 0.455 0.98 0.455 0.585 0.28 0.585 0.28 0.62 0.215 0.62  ;
  END
END CLKBUFX1

MACRO BUFX1  #BUF_X1
  CLASS core ;
  #FOREIGN BUF_X1 0.0 0.0 ;
  FOREIGN BUFX1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN Y  #Z
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.845 0.085 0.845 0.085 0.54 0.045 0.54 0.045 0.44 0.05 0.44 0.05 0.305 0.115 0.305 0.115 0.34 0.15 0.34 0.15 0.945 0.115 0.945 0.115 0.98 0.05 0.98  ;
    END
  END Y  #Z
  PIN A
    DIRECTION INPUT ;
	CAPACITANCE 0.000669 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.255 0.685 0.39 0.685 0.39 0.82 0.255 0.82  ;
    END
  END A
  PIN POWR #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 0.905 0.3 0.905 0.3 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.3 0.085 0.3 0.42 0.235 0.42 0.235 0.085 0 0.085  ;
    END
  END GRND  #VSS
  OBS
      LAYER M1 ;
        POLYGON 0.215 0.485 0.28 0.485 0.28 0.52 0.455 0.52 0.455 0.305 0.52 0.305 0.52 0.98 0.455 0.98 0.455 0.585 0.28 0.585 0.28 0.62 0.215 0.62  ;
  END
END BUFX1  #BUF_X1

MACRO BUFX2  #BUF_X2
  CLASS core ;
  #FOREIGN BUF_X2 0.0 0.0 ;
  FOREIGN BUFX2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN Y  #Z
    DIRECTION OUTPUT ;
	CAPACITANCE 0.016000 ;
    RESISTANCE 120.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.845 0.085 0.845 0.085 0.68 0.045 0.68 0.045 0.58 0.085 0.58 0.085 0.46 0.05 0.46 0.05 0.325 0.115 0.325 0.115 0.36 0.15 0.36 0.15 0.98 0.115 0.98 0.115 1.12 0.05 1.12  ;
    END
  END Y  #Z
  PIN A
    DIRECTION INPUT ;
	CAPACITANCE  0.000553 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.255 0.685 0.39 0.685 0.39 0.82 0.255 0.82  ;
    END
  END A
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 0.9 0.3 0.9 0.3 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.3 0.085 0.3 0.355 0.235 0.355 0.235 0.085 0 0.085  ;
    END
  END GRND  #VSS
  OBS
      LAYER M1 ;
        POLYGON 0.215 0.485 0.28 0.485 0.28 0.52 0.455 0.52 0.455 0.325 0.52 0.325 0.52 0.98 0.455 0.98 0.455 0.585 0.28 0.585 0.28 0.62 0.215 0.62  ;
  END
END BUFX2  #BUF_X2

MACRO BUFX3
  CLASS core ;
  FOREIGN BUFX3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN Y  #Z
    DIRECTION OUTPUT ;
	CAPACITANCE 0.024000 ;
    RESISTANCE 80.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.045 0.58 0.05 0.58 0.05 0.55 0.05 0.275 0.115 0.275 0.115 0.415 0.15 0.415 0.15 0.87 0.115 0.87 0.115 1.01 0.05 1.01 0.05 0.735 0.05 0.68 0.045 0.68  ;
    END
  END Y  #Z
  PIN A
    DIRECTION INPUT ;
	CAPACITANCE  0.000500 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.39 0.965 0.525 0.965 0.525 1.1 0.39 1.1  ;
    END
  END A
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 1.06 0.3 1.06 0.3 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.3 0.085 0.3 0.405 0.235 0.405 0.235 0.085 0 0.085  ;
    END
  END GRND  #VSS
  OBS
      LAYER M1 ;
        POLYGON 0.215 0.575 0.28 0.575 0.28 0.61 0.455 0.61 0.455 0.415 0.52 0.415 0.52 0.87 0.455 0.87 0.455 0.675 0.28 0.675 0.28 0.71 0.215 0.71  ;
  END
END BUFX3

MACRO BUFX4  #BUF_X4
  CLASS core ;
  #FOREIGN BUF_X4 0.0 0.0 ;
  FOREIGN BUFX4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN Y  #Z
    DIRECTION OUTPUT ;
	CAPACITANCE 0.032000 ;
    RESISTANCE 60.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.045 0.58 0.05 0.58 0.05 0.55 0.05 0.275 0.115 0.275 0.115 0.415 0.15 0.415 0.15 0.87 0.115 0.87 0.115 1.01 0.05 1.01 0.05 0.735 0.05 0.68 0.045 0.68  ;
    END
  END Y  #Z
  PIN A
    DIRECTION INPUT ;
	CAPACITANCE  0.000434 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.39 0.965 0.525 0.965 0.525 1.1 0.39 1.1  ;
    END
  END A
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 1.06 0.3 1.06 0.3 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.3 0.085 0.3 0.405 0.235 0.405 0.235 0.085 0 0.085  ;
    END
  END GRND  #VSS
  OBS
      LAYER M1 ;
        POLYGON 0.215 0.575 0.28 0.575 0.28 0.61 0.455 0.61 0.455 0.415 0.52 0.415 0.52 0.87 0.455 0.87 0.455 0.675 0.28 0.675 0.28 0.71 0.215 0.71  ;
  END
END BUFX4  #BUF_X4

MACRO BUFX8  #BUF_X8
  CLASS core ;
  #FOREIGN BUF_X8 0.0 0.0 ;
  FOREIGN BUFX8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN Y  #Z
    DIRECTION OUTPUT ;
	CAPACITANCE 0.064000 ;
    RESISTANCE 30.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.455 0.86 0.51 0.86 0.51 0.495 0.455 0.495 0.455 0.22 0.52 0.22 0.52 0.43 0.575 0.43 0.575 0.925 0.52 0.925 0.52 1.135 0.455 1.135  ;
    END
  END Y  #Z
  PIN A
    DIRECTION INPUT ;
	CAPACITANCE 0.001056 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.18 0.545 0.28 0.545 0.28 0.68 0.18 0.68  ;
    END
  END A
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.265 1.315 0.265 1.045 0.33 1.045 0.33 1.315 0.64 1.315 0.64 1.045 0.705 1.045 0.705 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.705 0.085 0.705 0.39 0.64 0.39 0.64 0.085 0.33 0.085 0.33 0.39 0.265 0.39 0.265 0.085 0 0.085  ;
    END
  END GRND  #VSS
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.385 0.115 0.385 0.115 0.745 0.345 0.745 0.345 0.595 0.38 0.595 0.38 0.56 0.445 0.56 0.445 0.695 0.41 0.695 0.41 0.81 0.115 0.81 0.115 0.88 0.05 0.88  ;
  END
END BUFX8  #BUF_X8

MACRO BUFX16  #BUF_X16
  CLASS core ;
  #FOREIGN BUF_X16 0.0 0.0 ;
  FOREIGN BUFX16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN Y  #Z
    DIRECTION OUTPUT ;
	CAPACITANCE 0.128000 ;
    RESISTANCE 15.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.445 0.275 0.51 0.275 0.51 0.485 0.82 0.485 0.82 0.275 0.885 0.275 0.885 0.58 0.905 0.58 0.905 0.68 0.885 0.68 0.885 1.01 0.82 1.01 0.82 0.68 0.805 0.68 0.805 0.58 0.805 0.55 0.51 0.55 0.51 1.01 0.445 1.01  ;
    END
  END Y  #Z
  PIN A
    DIRECTION INPUT ;
	CAPACITANCE 0.000412 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.06 0.965 0.16 0.965 0.16 1.1 0.06 1.1  ;
    END
  END A
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.255 1.315 0.255 1.06 0.32 1.06 0.32 1.315 0.635 1.315 0.635 1.06 0.7 1.06 0.7 1.315 1.01 1.315 1.01 1.06 1.075 1.06 1.075 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 1.075 0.085 1.075 0.405 1.01 0.405 1.01 0.085 0.695 0.085 0.695 0.405 0.63 0.405 0.63 0.085 0.32 0.085 0.32 0.405 0.255 0.405 0.255 0.085 0 0.085  ;
    END
  END GRND  #VSS
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.415 0.115 0.415 0.115 0.61 0.315 0.61 0.315 0.575 0.38 0.575 0.38 0.71 0.315 0.71 0.315 0.675 0.115 0.675 0.115 0.87 0.05 0.87  ;
  END
END BUFX16  #BUF_X16

MACRO BUFX32  #BUF_X32
  CLASS core ;
  #FOREIGN BUF_X32 0.0 0.0 ;
  FOREIGN BUFX32 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.9 BY 1.4 ;
  PIN Y  #Z
    DIRECTION OUTPUT ;
	CAPACITANCE 0.256000 ;
    RESISTANCE 7.5 ;
    PORT
      LAYER M1 ;
        POLYGON 0.715 0.58 0.715 0.645 1.785 0.645 1.785 0.92 1.72 0.92 1.72 0.71 1.405 0.71 1.405 0.92 1.34 0.92 1.34 0.71 1.025 0.71 1.025 0.92 0.96 0.92 0.96 0.71 0.65 0.71 0.65 0.92 0.585 0.92 0.585 0.28 0.65 0.28 0.65 0.49 0.96 0.49 0.96 0.28 1.025 0.28 1.025 0.49 1.34 0.49 1.34 0.28 1.405 0.28 1.405 0.49 1.72 0.49 1.72 0.28 1.785 0.28 1.785 0.555 0.715 0.555  ;
    END
  END Y  #Z
  PIN A
    DIRECTION INPUT ;
	CAPACITANCE 0.000434 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.27 0.31 0.37 0.31 0.37 1.09 0.27 1.09  ;
    END
  END A
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.395 1.315 0.395 1.185 0.46 1.185 0.46 1.315 0.77 1.315 0.77 1.045 0.835 1.045 0.835 1.315 1.15 1.315 1.15 1.045 1.215 1.045 1.215 1.315 1.53 1.315 1.53 1.045 1.595 1.045 1.595 1.315 1.9 1.315 1.9 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.9 -0.085 1.9 0.085 1.595 0.085 1.595 0.36 1.53 0.36 1.53 0.085 1.215 0.085 1.215 0.36 1.15 0.36 1.15 0.085 0.835 0.085 0.835 0.36 0.77 0.36 0.77 0.085 0.46 0.085 0.46 0.22 0.395 0.22 0.395 0.085 0 0.085  ;
    END
  END GRND  #VSS
  OBS
      LAYER M1 ;
        POLYGON 0.115 1.115 0.21 1.115 0.21 1.25 0.145 1.25 0.145 1.215 0.05 1.215 0.05 0.185 0.145 0.185 0.145 0.15 0.21 0.15 0.21 0.285 0.115 0.285  ;
  END
END BUFX32  #BUF_X32

MACRO OAI222_X1
  CLASS core ;
  FOREIGN OAI222_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.425 1.315 0.425 1.155 0.49 1.155 0.49 1.315 1.325 1.315 1.325 1.155 1.39 1.155 1.39 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.895 0.44 0.995 0.44 0.995 0.575 0.895 0.575  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.98 0.685 1.08 0.685 1.08 0.82 0.98 0.82  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.275 0.58 1.41 0.58 1.41 0.715 1.275 0.715  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 1.025 1.145 1.025 1.145 0.28 1.21 0.28 1.21 0.86 1.285 0.86 1.285 0.96 1.21 0.96 1.21 1.09 1.01 1.09 1.01 1.165 0.945 1.165 0.945 1.09 0.115 1.09 0.115 1.165 0.05 1.165  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.095 0.685 0.195 0.685 0.195 0.82 0.095 0.82  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 0.49 0.085 0.49 0.385 0.425 0.385 0.425 0.085 0.115 0.085 0.115 0.385 0.05 0.385 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.615 0.825 0.715 0.825 0.715 0.96 0.615 0.96  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.285 0.58 0.385 0.58 0.385 0.715 0.285 0.715  ;
    END
  END C2
  OBS
      LAYER M1 ;
        POLYGON 0.24 0.345 0.305 0.345 0.305 0.45 0.765 0.45 0.765 0.28 0.83 0.28 0.83 0.515 0.24 0.515  ;
        POLYGON 0.58 0.15 1.4 0.15 1.4 0.32 1.335 0.32 1.335 0.215 1.02 0.215 1.02 0.32 0.955 0.32 0.955 0.215 0.645 0.215 0.645 0.32 0.58 0.32  ;
  END
END OAI222_X1

MACRO OAI222_X2
  CLASS core ;
  FOREIGN OAI222_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.425 1.315 0.425 1.025 0.49 1.025 0.49 1.315 1.325 1.315 1.325 1.025 1.39 1.025 1.39 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.805 0.685 0.905 0.685 0.905 0.82 0.805 0.82  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.98 0.685 1.08 0.685 1.08 0.82 0.98 0.82  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.275 0.58 1.375 0.58 1.375 0.715 1.275 0.715  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.885 1.145 0.885 1.145 0.28 1.21 0.28 1.21 0.95 1.095 0.95 1.095 1 1.095 1.1 1.01 1.1 1.01 1.16 0.945 1.16 0.945 0.95 0.115 0.95 0.115 1.16 0.05 1.16  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.075 0.58 0.175 0.58 0.175 0.715 0.075 0.715  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 0.49 0.085 0.49 0.43 0.425 0.43 0.425 0.085 0.115 0.085 0.115 0.43 0.05 0.43 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.615 0.685 0.715 0.685 0.715 0.82 0.615 0.82  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.285 0.685 0.385 0.685 0.385 0.82 0.285 0.82  ;
    END
  END C2
  OBS
      LAYER M1 ;
        POLYGON 0.24 0.28 0.305 0.28 0.305 0.495 0.765 0.495 0.765 0.28 0.83 0.28 0.83 0.56 0.24 0.56  ;
        POLYGON 0.58 0.15 1.4 0.15 1.4 0.43 1.335 0.43 1.335 0.215 1.02 0.215 1.02 0.43 0.955 0.43 0.955 0.215 0.645 0.215 0.645 0.43 0.58 0.43  ;
  END
END OAI222_X2

MACRO OAI222_X4
  CLASS core ;
  FOREIGN OAI222_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 2.09 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.49 1.315 0.49 1.155 0.555 1.155 0.555 1.315 1.36 1.315 1.36 1.155 1.425 1.155 1.425 1.315 1.775 1.315 1.775 1.06 1.84 1.06 1.84 1.315 2.09 1.315 2.09 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.84 0.825 0.94 0.825 0.94 0.96 0.84 0.96  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.975 0.44 1.11 0.44 1.11 0.575 0.975 0.575  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.305 0.545 1.405 0.545 1.405 0.68 1.305 0.68  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.925 0.415 1.96 0.415 1.96 0.275 2.025 0.275 2.025 0.58 2.045 0.58 2.045 0.68 2.025 0.68 2.025 1.01 1.96 1.01 1.96 0.87 1.925 0.87  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.075 0.44 0.175 0.44 0.175 0.575 0.075 0.575  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 2.09 -0.085 2.09 0.085 1.84 0.085 1.84 0.405 1.775 0.405 1.775 0.085 0.49 0.085 0.49 0.32 0.425 0.32 0.425 0.085 0.115 0.085 0.115 0.32 0.05 0.32 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.615 0.685 0.715 0.685 0.715 0.82 0.615 0.82  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.35 0.545 0.45 0.545 0.45 0.68 0.35 0.68  ;
    END
  END C2
  OBS
      LAYER M1 ;
        POLYGON 0.24 0.28 0.305 0.28 0.305 0.385 0.765 0.385 0.765 0.28 0.83 0.28 0.83 0.45 0.24 0.45  ;
        POLYGON 0.58 0.15 1.425 0.15 1.425 0.32 1.36 0.32 1.36 0.215 1.02 0.215 1.02 0.32 0.955 0.32 0.955 0.215 0.645 0.215 0.645 0.32 0.58 0.32  ;
        POLYGON 0.115 1.025 1.175 1.025 1.175 0.28 1.24 0.28 1.24 0.745 1.465 0.745 1.465 0.71 1.53 0.71 1.53 0.845 1.465 0.845 1.465 0.81 1.24 0.81 1.24 1.09 1.025 1.09 1.025 1.165 0.96 1.165 0.96 1.09 0.18 1.09 0.18 1.165 0.115 1.165  ;
        POLYGON 1.555 0.905 1.595 0.905 1.595 0.55 1.555 0.55 1.555 0.415 1.62 0.415 1.62 0.49 1.66 0.49 1.66 0.61 1.795 0.61 1.795 0.575 1.86 0.575 1.86 0.71 1.795 0.71 1.795 0.675 1.66 0.675 1.66 0.965 1.62 0.965 1.62 1.18 1.555 1.18  ;
  END
END OAI222_X4

MACRO AND3_X1
  CLASS core ;
  FOREIGN AND3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.25 1.315 0.25 1.07 0.315 1.07 0.315 1.315 0.645 1.315 0.645 1.07 0.71 1.07 0.71 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.34 0.44 0.44 0.44 0.44 0.575 0.34 0.575  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.67 0.685 0.77 0.685 0.77 0.82 0.67 0.82  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.335 0.085 0.335 0.32 0.27 0.32 0.27 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.505 0.545 0.605 0.545 0.605 0.68 0.505 0.68  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 1.01 0.085 1.01 0.085 0.54 0.045 0.54 0.045 0.44 0.05 0.44 0.05 0.415 0.05 0.28 0.115 0.28 0.115 0.315 0.15 0.315 0.15 1.11 0.115 1.11 0.115 1.145 0.05 1.145  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.215 0.85 0.28 0.85 0.28 0.885 0.835 0.885 0.835 0.28 0.9 0.28 0.9 1.145 0.835 1.145 0.835 0.95 0.525 0.95 0.525 1.145 0.46 1.145 0.46 0.95 0.28 0.95 0.28 0.985 0.215 0.985  ;
  END
END AND3_X1

MACRO AND3_X2
  CLASS core ;
  FOREIGN AND3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 0.925 0.3 0.925 0.3 1.315 0.645 1.315 0.645 0.93 0.71 0.93 0.71 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.315 0.44 0.415 0.44 0.415 0.575 0.315 0.575  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.67 0.44 0.77 0.44 0.77 0.575 0.67 0.575  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.3 0.085 0.3 0.31 0.235 0.31 0.235 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.505 0.545 0.605 0.545 0.605 0.68 0.505 0.68  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.87 0.085 0.87 0.085 0.54 0.045 0.54 0.045 0.44 0.05 0.44 0.05 0.415 0.05 0.28 0.115 0.28 0.115 0.315 0.15 0.315 0.15 1.005 0.115 1.005 0.115 1.145 0.05 1.145  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.215 0.71 0.28 0.71 0.28 0.745 0.835 0.745 0.835 0.28 0.9 0.28 0.9 1.005 0.835 1.005 0.835 0.81 0.525 0.81 0.525 1.005 0.46 1.005 0.46 0.81 0.28 0.81 0.28 0.845 0.215 0.845  ;
  END
END AND3_X2

MACRO AND3_X4
  CLASS core ;
  FOREIGN AND3_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 1.06 0.3 1.06 0.3 1.315 0.645 1.315 0.645 1.015 0.71 1.015 0.71 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.375 0.405 0.475 0.405 0.475 0.54 0.375 0.54  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.67 0.545 0.77 0.545 0.77 0.68 0.67 0.68  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.3 0.085 0.3 0.265 0.235 0.265 0.235 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.505 0.685 0.605 0.685 0.605 0.82 0.505 0.82  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.045 0.58 0.05 0.58 0.05 0.55 0.05 0.275 0.115 0.275 0.115 0.415 0.15 0.415 0.15 0.87 0.115 0.87 0.115 1.01 0.05 1.01 0.05 0.735 0.05 0.68 0.045 0.68  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.215 0.575 0.28 0.575 0.28 0.885 0.835 0.885 0.835 0.225 0.9 0.225 0.9 1.09 0.835 1.09 0.835 0.95 0.525 0.95 0.525 1.09 0.46 1.09 0.46 0.95 0.215 0.95  ;
  END
END AND3_X4

MACRO AOI221_X1
  CLASS core ;
  FOREIGN AOI221_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.445 0.67 0.58 0.67 0.58 0.805 0.445 0.805  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.83 1.315 0.83 0.875 0.895 0.875 0.895 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.715 0.545 0.815 0.545 0.815 0.68 0.715 0.68  ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.165 0.115 0.165 0.115 0.31 0.64 0.31 0.64 0.165 0.705 0.165 0.705 0.375 0.3 0.375 0.3 0.72 0.335 0.72 0.335 0.82 0.3 0.82 0.3 1.105 0.235 1.105 0.235 0.82 0.235 0.72 0.235 0.375 0.05 0.375  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.07 0.58 0.17 0.58 0.17 0.715 0.07 0.715  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 1.085 0.085 1.085 0.245 1.02 0.245 1.02 0.085 0.49 0.085 0.49 0.245 0.425 0.245 0.425 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.88 0.405 0.98 0.405 0.98 0.54 0.88 0.54  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.44 0.5 0.44 0.5 0.575 0.365 0.575  ;
    END
  END C2
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.875 0.115 0.875 0.115 1.17 0.425 1.17 0.425 0.875 0.49 0.875 0.49 1.235 0.05 1.235  ;
        POLYGON 0.645 0.745 1.085 0.745 1.085 1.105 1.02 1.105 1.02 0.81 0.71 0.81 0.71 1.105 0.645 1.105  ;
  END
END AOI221_X1

MACRO AOI221_X2
  CLASS core ;
  FOREIGN AOI221_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.58 0.665 0.58 0.665 0.68 0.53 0.68  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.82 1.315 0.82 1.035 0.885 1.035 0.885 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.73 0.57 0.83 0.57 0.83 0.705 0.73 0.705  ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.255 0.115 0.255 0.115 0.41 0.63 0.41 0.63 0.255 0.695 0.255 0.695 0.475 0.3 0.475 0.3 0.86 0.335 0.86 0.335 0.96 0.3 0.96 0.3 1.005 0.235 1.005 0.235 0.96 0.235 0.86 0.235 0.475 0.05 0.475  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.07 0.57 0.17 0.57 0.17 0.705 0.07 0.705  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 1.075 0.085 1.075 0.345 1.01 0.345 1.01 0.085 0.49 0.085 0.49 0.345 0.425 0.345 0.425 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.87 0.415 1.005 0.415 1.005 0.515 0.87 0.515  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.57 0.465 0.57 0.465 0.705 0.365 0.705  ;
    END
  END C2
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.86 0.115 0.86 0.115 1.07 0.425 1.07 0.425 0.86 0.49 0.86 0.49 1.135 0.05 1.135  ;
        POLYGON 0.635 0.905 1.075 0.905 1.075 1.04 1.01 1.04 1.01 0.97 0.7 0.97 0.7 1.04 0.635 1.04  ;
  END
END AOI221_X2

MACRO AOI221_X4
  CLASS core ;
  FOREIGN AOI221_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.71 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.495 0.44 0.595 0.44 0.595 0.575 0.495 0.575  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.84 1.315 0.84 0.885 0.905 0.885 0.905 1.315 1.405 1.315 1.405 1.055 1.47 1.055 1.47 1.315 1.71 1.315 1.71 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.79 0.405 0.89 0.405 0.89 0.54 0.79 0.54  ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.555 0.41 1.59 0.41 1.59 0.27 1.655 0.27 1.655 0.58 1.665 0.58 1.665 0.68 1.655 0.68 1.655 1.005 1.59 1.005 1.59 0.865 1.555 0.865  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.07 0.58 0.17 0.58 0.17 0.715 0.07 0.715  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.71 -0.085 1.71 0.085 1.47 0.085 1.47 0.4 1.405 0.4 1.405 0.085 1.1 0.085 1.1 0.28 1.035 0.28 1.035 0.085 0.49 0.085 0.49 0.245 0.425 0.245 0.425 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.955 0.405 1.055 0.405 1.055 0.54 0.955 0.54  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.64 0.5 0.64 0.5 0.775 0.365 0.775  ;
    END
  END C2
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.885 0.115 0.885 0.115 1.18 0.425 1.18 0.425 0.885 0.49 0.885 0.49 1.245 0.05 1.245  ;
        POLYGON 0.655 0.755 1.095 0.755 1.095 1.115 1.03 1.115 1.03 0.82 0.72 0.82 0.72 1.115 0.655 1.115  ;
        POLYGON 0.05 0.165 0.115 0.165 0.115 0.31 0.66 0.31 0.66 0.2 0.725 0.2 0.725 0.605 1.14 0.605 1.14 0.57 1.205 0.57 1.205 0.705 1.14 0.705 1.14 0.67 0.66 0.67 0.66 0.375 0.3 0.375 0.3 1.115 0.235 1.115 0.235 0.375 0.05 0.375  ;
        POLYGON 1.185 0.77 1.27 0.77 1.27 0.505 1.185 0.505 1.185 0.37 1.25 0.37 1.25 0.405 1.335 0.405 1.335 0.605 1.425 0.605 1.425 0.57 1.49 0.57 1.49 0.705 1.425 0.705 1.425 0.67 1.335 0.67 1.335 0.905 1.25 0.905 1.25 1.045 1.185 1.045  ;
  END
END AOI221_X4

MACRO NOR4X1  #NOR4_X1
  CLASS core ;
  #FOREIGN NOR4_X1 0.0 0.0 ;
  FOREIGN NOR4X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.805 1.315 0.805 0.955 0.87 0.955 0.87 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN C  #A3
    DIRECTION INPUT ;
	CAPACITANCE 0.000373 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.5 0.545 0.6 0.545 0.6 0.68 0.5 0.68  ;
    END
  END C  #A3
  PIN A  #A1
    DIRECTION INPUT ;
	CAPACITANCE 0.000389 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.18 0.685 0.28 0.685 0.28 0.82 0.18 0.82  ;
    END
  END A  #A1
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.87 0.085 0.87 0.29 0.805 0.29 0.805 0.085 0.49 0.085 0.49 0.29 0.425 0.29 0.425 0.085 0.115 0.085 0.115 0.29 0.05 0.29 0.05 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN B  #A2
    DIRECTION INPUT ;
	CAPACITANCE 0.000669 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.285 0.485 0.385 0.485 0.385 0.62 0.285 0.62  ;
    END
  END B  #A2
  PIN D  #A4
    DIRECTION INPUT ;
	CAPACITANCE 0.000360 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.665 0.685 0.765 0.685 0.765 0.82 0.665 0.82  ;
    END
  END D  #A4
  PIN Y  #ZN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.355 0.24 0.355 0.24 0.175 0.305 0.175 0.305 0.355 0.615 0.355 0.615 0.26 0.615 0.175 0.615 0.16 0.715 0.16 0.715 0.26 0.68 0.26 0.68 0.42 0.115 0.42 0.115 1.12 0.05 1.12  ;
    END
  END Y  #ZN
END NOR4X1  #NOR4_X1

MACRO NOR4_X2
  CLASS core ;
  FOREIGN NOR4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.805 1.315 0.805 1.06 0.87 1.06 0.87 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.51 0.44 0.61 0.44 0.61 0.575 0.51 0.575  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.18 0.44 0.28 0.44 0.28 0.575 0.18 0.575  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.87 0.085 0.87 0.245 0.805 0.245 0.805 0.085 0.49 0.085 0.49 0.245 0.425 0.245 0.425 0.085 0.115 0.085 0.115 0.245 0.05 0.245 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.345 0.44 0.445 0.44 0.445 0.575 0.345 0.575  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.725 0.44 0.825 0.44 0.825 0.575 0.725 0.575  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.31 0.24 0.31 0.24 0.215 0.305 0.215 0.305 0.31 0.615 0.31 0.615 0.215 0.68 0.215 0.68 0.375 0.115 0.375 0.115 0.9 0.05 0.9  ;
    END
  END ZN
END NOR4_X2

MACRO NOR4_X4
  CLASS core ;
  FOREIGN NOR4_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.71 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.04 1.315 0.04 1.095 0.175 1.095 0.175 1.315 1.59 1.315 1.59 1.06 1.655 1.06 1.655 1.315 1.71 1.315 1.71 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.465 0.435 0.465 0.435 0.705 1.295 0.705 1.295 0.465 1.36 0.465 1.36 0.77 0.37 0.77  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.77 0.375 0.905 0.375 0.905 0.51 0.77 0.51  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.71 -0.085 1.71 0.085 1.655 0.085 1.655 0.215 1.59 0.215 1.59 0.085 1.31 0.085 1.31 0.18 1.175 0.18 1.175 0.085 0.93 0.085 0.93 0.18 0.795 0.18 0.795 0.085 0.55 0.085 0.55 0.18 0.415 0.18 0.415 0.085 0.175 0.085 0.175 0.18 0.04 0.18 0.04 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.56 0.465 0.625 0.465 0.625 0.575 1.105 0.575 1.105 0.465 1.17 0.465 1.17 0.64 0.56 0.64  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.21 0.465 0.275 0.465 0.275 0.835 1.485 0.835 1.485 0.465 1.55 0.465 1.55 0.9 1.095 0.9 1.095 0.96 0.995 0.96 0.995 0.9 0.21 0.9  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.045 0.44 0.08 0.44 0.08 0.245 0.265 0.245 0.265 0.175 0.33 0.175 0.33 0.245 0.645 0.245 0.645 0.175 0.71 0.175 0.71 0.245 1.025 0.245 1.025 0.175 1.09 0.175 1.09 0.245 1.4 0.245 1.4 0.175 1.465 0.175 1.465 0.31 0.145 0.31 0.145 0.44 0.145 0.54 0.145 0.965 0.895 0.965 0.895 1 0.93 1 0.93 1.205 0.795 1.205 0.795 1.03 0.08 1.03 0.08 0.54 0.045 0.54  ;
    END
  END ZN
END NOR4_X4

MACRO OAI211_X1
  CLASS core ;
  FOREIGN OAI211_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.535 0.55 0.635 0.55 0.635 0.685 0.535 0.685  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.11 0.115 1.11 0.115 1.315 0.63 1.315 0.63 1.11 0.695 1.11 0.695 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.87 0.085 0.87 0.32 0.805 0.32 0.805 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.69 0.72 0.825 0.72 0.825 0.855 0.69 0.855  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 1 0.24 1 0.24 0.28 0.305 0.28 0.305 0.98 0.895 0.98 0.895 1.185 0.83 1.185 0.83 1.045 0.49 1.045 0.49 1.12 0.425 1.12 0.425 1.045 0.335 1.045 0.335 1.1 0.235 1.1  ;
    END
  END ZN
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.075 0.825 0.175 0.825 0.175 0.96 0.075 0.96  ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.44 0.47 0.44 0.47 0.575 0.37 0.575  ;
    END
  END C1
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.15 0.49 0.15 0.49 0.32 0.425 0.32 0.425 0.215 0.115 0.215 0.115 0.32 0.05 0.32  ;
  END
END OAI211_X1

MACRO OAI211_X2
  CLASS core ;
  FOREIGN OAI211_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.545 0.685 0.645 0.685 0.645 0.82 0.545 0.82  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.025 0.115 1.025 0.115 1.315 0.63 1.315 0.63 1.015 0.695 1.015 0.695 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.885 0.085 0.885 0.43 0.82 0.43 0.82 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.71 0.58 0.81 0.58 0.81 0.715 0.71 0.715  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.25 0.28 0.315 0.28 0.315 0.885 0.885 0.885 0.885 1.235 0.82 1.235 0.82 0.95 0.525 0.95 0.525 1 0.525 1.1 0.49 1.1 0.49 1.16 0.425 1.16 0.425 1.1 0.425 1 0.425 0.95 0.25 0.95  ;
    END
  END ZN
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.085 0.685 0.185 0.685 0.185 0.82 0.085 0.82  ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.38 0.58 0.48 0.58 0.48 0.715 0.38 0.715  ;
    END
  END C1
  OBS
      LAYER M1 ;
        POLYGON 0.065 0.15 0.505 0.15 0.505 0.43 0.44 0.43 0.44 0.215 0.13 0.215 0.13 0.43 0.065 0.43  ;
  END
END OAI211_X2

MACRO OAI211_X4
  CLASS core ;
  FOREIGN OAI211_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.515 0.825 0.615 0.825 0.615 0.96 0.515 0.96  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.155 0.115 1.155 0.115 1.315 0.63 1.315 0.63 1.155 0.695 1.155 0.695 1.315 1.22 1.315 1.22 1.06 1.285 1.06 1.285 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 1.285 0.085 1.285 0.405 1.22 0.405 1.22 0.085 0.885 0.085 0.885 0.32 0.82 0.32 0.82 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.68 0.44 0.815 0.44 0.815 0.575 0.68 0.575  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.37 0.415 1.405 0.415 1.405 0.275 1.47 0.275 1.47 0.58 1.475 0.58 1.475 0.68 1.47 0.68 1.47 1.01 1.405 1.01 1.405 0.87 1.37 0.87  ;
    END
  END ZN
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.09 0.72 0.19 0.72 0.19 0.855 0.09 0.855  ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.385 0.545 0.485 0.545 0.485 0.68 0.385 0.68  ;
    END
  END C1
  OBS
      LAYER M1 ;
        POLYGON 0.065 0.15 0.505 0.15 0.505 0.32 0.44 0.32 0.44 0.215 0.13 0.215 0.13 0.32 0.065 0.32  ;
        POLYGON 0.255 0.28 0.32 0.28 0.32 1.025 0.87 1.025 0.87 0.61 0.905 0.61 0.905 0.575 0.97 0.575 0.97 0.71 0.935 0.71 0.935 1.23 0.82 1.23 0.82 1.09 0.49 1.09 0.49 1.165 0.425 1.165 0.425 1.09 0.255 1.09  ;
        POLYGON 1 0.77 1.035 0.77 1.035 0.515 1 0.515 1 0.38 1.065 0.38 1.065 0.415 1.1 0.415 1.1 0.61 1.24 0.61 1.24 0.575 1.305 0.575 1.305 0.71 1.24 0.71 1.24 0.675 1.1 0.675 1.1 0.905 1.065 0.905 1.065 1.045 1 1.045  ;
  END
END OAI211_X4

MACRO AND4_X1
  CLASS core ;
  FOREIGN AND4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.25 1.315 0.25 1.155 0.315 1.155 0.315 1.315 0.645 1.315 0.645 1.155 0.71 1.155 0.71 1.315 1.025 1.315 1.025 1.155 1.09 1.155 1.09 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.505 0.825 0.605 0.825 0.605 0.96 0.505 0.96  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.86 0.685 0.96 0.685 0.96 0.82 0.86 0.82  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.335 0.085 0.335 0.275 0.27 0.275 0.27 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.695 0.545 0.795 0.545 0.795 0.68 0.695 0.68  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.315 0.44 0.415 0.44 0.415 0.575 0.315 0.575  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 1.095 0.085 1.095 0.085 0.54 0.045 0.54 0.045 0.44 0.05 0.44 0.05 0.415 0.05 0.28 0.115 0.28 0.115 0.315 0.15 0.315 0.15 1.195 0.115 1.195 0.115 1.23 0.05 1.23  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.215 0.935 0.28 0.935 0.28 1.025 1.025 1.025 1.025 0.28 1.09 0.28 1.09 1.09 0.905 1.09 0.905 1.23 0.84 1.23 0.84 1.09 0.525 1.09 0.525 1.23 0.46 1.23 0.46 1.09 0.215 1.09  ;
  END
END AND4_X1

MACRO AND4_X2
  CLASS core ;
  FOREIGN AND4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 1.015 0.3 1.015 0.3 1.315 0.645 1.315 0.645 1.02 0.71 1.02 0.71 1.315 1.025 1.315 1.025 1.02 1.09 1.02 1.09 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.505 0.685 0.605 0.685 0.605 0.82 0.505 0.82  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.86 0.545 0.96 0.545 0.96 0.68 0.86 0.68  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.335 0.085 0.335 0.275 0.27 0.275 0.27 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.695 0.44 0.795 0.44 0.795 0.575 0.695 0.575  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.315 0.58 0.415 0.58 0.415 0.715 0.315 0.715  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.96 0.085 0.96 0.085 0.54 0.045 0.54 0.045 0.44 0.05 0.44 0.05 0.415 0.05 0.28 0.115 0.28 0.115 0.315 0.15 0.315 0.15 1.095 0.115 1.095 0.115 1.235 0.05 1.235  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.215 0.8 0.28 0.8 0.28 0.885 0.485 0.885 0.485 0.89 1.025 0.89 1.025 0.28 1.09 0.28 1.09 0.955 0.905 0.955 0.905 1.095 0.84 1.095 0.84 0.955 0.525 0.955 0.525 1.095 0.46 1.095 0.46 0.95 0.215 0.95  ;
  END
END AND4_X2

MACRO AND4_X4
  CLASS core ;
  FOREIGN AND4_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 1.045 0.3 1.045 0.3 1.315 0.645 1.315 0.645 1.015 0.71 1.015 0.71 1.315 1.025 1.315 1.025 1.015 1.09 1.015 1.09 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.505 0.685 0.605 0.685 0.605 0.82 0.505 0.82  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.86 0.685 0.96 0.685 0.96 0.82 0.86 0.82  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.3 0.085 0.3 0.39 0.235 0.39 0.235 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.72 0.44 0.82 0.44 0.82 0.575 0.72 0.575  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.345 0.44 0.445 0.44 0.445 0.575 0.345 0.575  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.045 0.58 0.05 0.58 0.05 0.535 0.05 0.26 0.115 0.26 0.115 0.4 0.15 0.4 0.15 0.855 0.115 0.855 0.115 0.995 0.05 0.995 0.05 0.72 0.05 0.68 0.045 0.68  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.215 0.56 0.28 0.56 0.28 0.885 1.025 0.885 1.025 0.28 1.09 0.28 1.09 0.95 0.905 0.95 0.905 1.09 0.84 1.09 0.84 0.95 0.525 0.95 0.525 1.09 0.46 1.09 0.46 0.95 0.215 0.95  ;
  END
END AND4_X4

MACRO NAND3X1  #NAND3_X1
  CLASS core ;
  #FOREIGN NAND3_X1 0.0 0.0 ;
  FOREIGN NAND3X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 1.015 0.3 1.015 0.3 1.315 0.615 1.315 0.615 1.015 0.68 1.015 0.68 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN C  #A3
    DIRECTION INPUT ;
	CAPACITANCE 0.000347 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.51 0.685 0.61 0.685 0.61 0.82 0.51 0.82  ;
    END
  END C  #A3
  PIN A  #A1
    DIRECTION INPUT ;
	CAPACITANCE 0.000390 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.18 0.44 0.28 0.44 0.28 0.575 0.18 0.575  ;
    END
  END A  #A1
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.68 0.085 0.68 0.32 0.615 0.32 0.615 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN B  #A2
    DIRECTION INPUT ;
	CAPACITANCE 0.000360 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.345 0.545 0.445 0.545 0.445 0.68 0.345 0.68  ;
    END
  END B  #A2
  PIN Y  #ZN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.28 0.115 0.28 0.115 0.885 0.49 0.885 0.49 1 0.525 1 0.525 1.1 0.425 1.1 0.425 1.09 0.425 1 0.425 0.95 0.115 0.95 0.115 1.09 0.05 1.09  ;
    END
  END Y  #ZN
END NAND3X1  #NAND3_X1

MACRO NAND3_X2
  CLASS core ;
  FOREIGN NAND3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 1.015 0.3 1.015 0.3 1.315 0.615 1.315 0.615 1.015 0.68 1.015 0.68 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.51 0.58 0.61 0.58 0.61 0.715 0.51 0.715  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.18 0.58 0.28 0.58 0.28 0.715 0.18 0.715  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.68 0.085 0.68 0.43 0.615 0.43 0.615 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.345 0.685 0.445 0.685 0.445 0.82 0.345 0.82  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.28 0.115 0.28 0.115 0.885 0.49 0.885 0.49 1 0.525 1 0.525 1.1 0.49 1.1 0.49 1.235 0.425 1.235 0.425 1.1 0.425 1 0.425 0.95 0.115 0.95 0.115 1.235 0.05 1.235  ;
    END
  END ZN
END NAND3_X2

MACRO NAND3_X4
  CLASS core ;
  FOREIGN NAND3_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.06 0.115 1.06 0.115 1.315 0.39 1.315 0.39 1.235 0.525 1.235 0.525 1.315 0.77 1.315 0.77 1.235 0.905 1.235 0.905 1.315 1.15 1.315 1.15 1.235 1.285 1.235 1.285 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.535 0.845 0.765 0.845 0.765 0.98 0.7 0.98 0.7 0.91 0.6 0.91 0.6 0.98 0.535 0.98  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.155 0.585 1.115 0.585 1.115 0.72 1.05 0.72 1.05 0.65 0.22 0.65 0.22 0.72 0.155 0.72  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 1.15 0.185 1.185 0.185 1.185 0.085 0.115 0.085 0.115 0.425 0.05 0.425 0.05 0.085 0 0.085 0 -0.085 1.33 -0.085 1.33 0.085 1.25 0.085 1.25 0.185 1.285 0.185 1.285 0.39 1.15 0.39  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.345 0.715 0.955 0.715 0.955 0.85 0.89 0.85 0.89 0.78 0.41 0.78 0.41 0.85 0.345 0.85  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 1.045 0.995 1.045 0.995 1 1.095 1 1.095 1.045 1.18 1.045 1.18 0.52 0.62 0.52 0.62 0.485 0.585 0.485 0.585 0.28 0.72 0.28 0.72 0.455 1.245 0.455 1.245 1.11 1.065 1.11 1.065 1.18 1 1.18 1 1.11 0.685 1.11 0.685 1.18 0.62 1.18 0.62 1.11 0.305 1.11 0.305 1.18 0.24 1.18  ;
    END
  END ZN
END NAND3_X4

MACRO OR4X1  #OR4_X1
  CLASS core ;
  #FOREIGN OR4_X1 0.0 0.0 ;
  FOREIGN OR4X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.27 1.315 0.27 0.955 0.335 0.955 0.335 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN C  #A3
    DIRECTION INPUT ;
	CAPACITANCE 0.000515 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.58 0.63 0.58 0.63 0.715 0.53 0.715  ;
    END
  END C  #A3
  PIN A  #A1
    DIRECTION INPUT ;
	CAPACITANCE 0.000624 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.86 0.58 0.96 0.58 0.96 0.715 0.86 0.715  ;
    END
  END A  #A1
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 1.09 0.085 1.09 0.35 1.025 0.35 1.025 0.085 0.71 0.085 0.71 0.35 0.645 0.35 0.645 0.085 0.315 0.085 0.315 0.35 0.25 0.35 0.25 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN B  #A2
    DIRECTION INPUT ;
	CAPACITANCE 0.000374 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.695 0.685 0.795 0.685 0.795 0.82 0.695 0.82  ;
    END
  END B  #A2
  PIN D  #A4
    DIRECTION INPUT ;
	CAPACITANCE 0.000364 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.315 0.685 0.415 0.685 0.415 0.82 0.315 0.82  ;
    END
  END D  #A4
  PIN Y  #ZN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.845 0.085 0.845 0.085 0.54 0.045 0.54 0.045 0.44 0.085 0.44 0.085 0.37 0.05 0.37 0.05 0.235 0.115 0.235 0.115 0.27 0.15 0.27 0.15 0.945 0.115 0.945 0.115 0.98 0.05 0.98  ;
    END
  END Y  #ZN
  OBS
      LAYER M1 ;
        POLYGON 0.215 0.415 0.28 0.415 0.28 0.45 0.455 0.45 0.455 0.235 0.52 0.235 0.52 0.45 0.835 0.45 0.835 0.235 0.9 0.235 0.9 0.45 1.09 0.45 1.09 1.12 1.025 1.12 1.025 0.515 0.28 0.515 0.28 0.55 0.215 0.55  ;
  END
END OR4X1  #OR4_X1

MACRO OR4_X2
  CLASS core ;
  FOREIGN OR4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.27 1.315 0.27 0.955 0.335 0.955 0.335 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.53 0.58 0.63 0.58 0.63 0.715 0.53 0.715  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.86 0.58 0.96 0.58 0.96 0.715 0.86 0.715  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 1.09 0.085 1.09 0.37 1.025 0.37 1.025 0.085 0.71 0.085 0.71 0.37 0.645 0.37 0.645 0.085 0.3 0.085 0.3 0.285 0.235 0.285 0.235 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.695 0.685 0.795 0.685 0.795 0.82 0.695 0.82  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.315 0.685 0.415 0.685 0.415 0.82 0.315 0.82  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.845 0.085 0.845 0.085 0.54 0.045 0.54 0.045 0.44 0.05 0.44 0.05 0.39 0.05 0.255 0.115 0.255 0.115 0.29 0.15 0.29 0.15 0.98 0.115 0.98 0.115 1.12 0.05 1.12  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.215 0.415 0.28 0.415 0.28 0.45 0.455 0.45 0.455 0.255 0.52 0.255 0.52 0.45 0.835 0.45 0.835 0.255 0.9 0.255 0.9 0.45 1.09 0.45 1.09 1.12 1.025 1.12 1.025 0.515 0.28 0.515 0.28 0.55 0.215 0.55  ;
  END
END OR4_X2

MACRO OR4_X4
  CLASS core ;
  FOREIGN OR4_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 1.045 0.3 1.045 0.3 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.54 0.7 0.64 0.7 0.64 0.835 0.54 0.835  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.945 0.685 1.045 0.685 1.045 0.82 0.945 0.82  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 1.09 0.085 1.09 0.49 1.025 0.49 1.025 0.085 0.71 0.085 0.71 0.49 0.645 0.49 0.645 0.085 0.3 0.085 0.3 0.365 0.235 0.365 0.235 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.72 0.7 0.82 0.7 0.82 0.835 0.72 0.835  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.375 0.7 0.475 0.7 0.475 0.835 0.375 0.835  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.045 0.58 0.085 0.58 0.085 0.51 0.05 0.51 0.05 0.235 0.115 0.235 0.115 0.375 0.15 0.375 0.15 0.855 0.115 0.855 0.115 0.995 0.05 0.995 0.05 0.72 0.05 0.68 0.045 0.68  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.28 0.915 0.42 0.915 0.42 0.955 1.025 0.955 1.025 0.885 1.09 0.885 1.09 1.16 1.025 1.16 1.025 1.02 0.36 1.02 0.36 0.98 0.215 0.98 0.215 0.535 0.28 0.535 0.28 0.57 0.455 0.57 0.455 0.375 0.52 0.375 0.52 0.57 0.835 0.57 0.835 0.375 0.9 0.375 0.9 0.635 0.28 0.635  ;
  END
END OR4_X4

MACRO OAI21X1  #OAI21_X1
  CLASS core ;
  #FOREIGN OAI21_X1 0.0 0.0 ;
  FOREIGN OAI21X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN A0  #A
    DIRECTION INPUT ;
	CAPACITANCE 0.000365 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.535 0.825 0.635 0.825 0.635 0.96 0.535 0.96  ;
    END
  END A0  #A
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.11 0.115 1.11 0.115 1.315 0.615 1.315 0.615 1.045 0.68 1.045 0.68 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END POWR  #VDD
  PIN A1  #B1
    DIRECTION INPUT ;
	CAPACITANCE 0.000365 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.685 0.47 0.685 0.47 0.82 0.37 0.82  ;
    END
  END A1  #B1
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.68 0.085 0.68 0.5 0.615 0.5 0.615 0.085 0 0.085  ;
    END
  END GRND  #VSS
  PIN B0  #B2
    DIRECTION INPUT ;
	CAPACITANCE 0.000442 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.075 0.58 0.175 0.58 0.175 0.715 0.075 0.715  ;
    END
  END B0  #B2
  PIN Y  #ZN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 1 0.24 1 0.24 0.42 0.305 0.42 0.305 1 0.335 1 0.335 1.01 0.49 1.01 0.49 1.145 0.425 1.145 0.425 1.075 0.335 1.075 0.335 1.1 0.235 1.1  ;
    END
  END Y  #ZN
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.29 0.49 0.29 0.49 0.5 0.425 0.5 0.425 0.355 0.115 0.355 0.115 0.5 0.05 0.5  ;
  END
END OAI21X1  #OAI21_X1

MACRO OAI21_X2
  CLASS core ;
  FOREIGN OAI21_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.535 0.685 0.635 0.685 0.635 0.82 0.535 0.82  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.025 0.115 1.025 0.115 1.315 0.615 1.315 0.615 0.9 0.68 0.9 0.68 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.37 0.58 0.47 0.58 0.47 0.715 0.37 0.715  ;
    END
  END B1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.68 0.085 0.68 0.51 0.615 0.51 0.615 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.075 0.685 0.175 0.685 0.175 0.82 0.075 0.82  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.24 0.28 0.305 0.28 0.305 0.87 0.49 0.87 0.49 1 0.525 1 0.525 1.1 0.49 1.1 0.49 1.145 0.425 1.145 0.425 1.1 0.425 1 0.425 0.935 0.24 0.935  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.15 0.49 0.15 0.49 0.51 0.425 0.51 0.425 0.215 0.115 0.215 0.115 0.51 0.05 0.51  ;
  END
END OAI21_X2

MACRO OAI21_X4
  CLASS core ;
  FOREIGN OAI21_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.535 0.44 0.635 0.44 0.635 0.575 0.535 0.575  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.155 0.115 1.155 0.115 1.315 0.64 1.315 0.64 1.155 0.705 1.155 0.705 1.315 1.015 1.315 1.015 1.06 1.08 1.06 1.08 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.365 0.825 0.5 0.825 0.5 0.96 0.365 0.96  ;
    END
  END B1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 1.08 0.085 1.08 0.405 1.015 0.405 1.015 0.085 0.705 0.085 0.705 0.36 0.64 0.36 0.64 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.07 0.72 0.17 0.72 0.17 0.855 0.07 0.855  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.165 0.415 1.2 0.415 1.2 0.275 1.265 0.275 1.265 0.58 1.285 0.58 1.285 0.68 1.265 0.68 1.265 1.01 1.2 1.01 1.2 0.87 1.165 0.87  ;
    END
  END ZN
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.15 0.49 0.15 0.49 0.36 0.425 0.36 0.425 0.215 0.115 0.215 0.115 0.36 0.05 0.36  ;
        POLYGON 0.235 0.28 0.3 0.28 0.3 1.025 0.565 1.025 0.565 0.645 0.7 0.645 0.7 0.575 0.765 0.575 0.765 0.71 0.63 0.71 0.63 1.09 0.49 1.09 0.49 1.165 0.425 1.165 0.425 1.09 0.235 1.09  ;
        POLYGON 0.795 0.77 0.83 0.77 0.83 0.515 0.795 0.515 0.795 0.38 0.86 0.38 0.86 0.415 0.895 0.415 0.895 0.61 1.035 0.61 1.035 0.575 1.1 0.575 1.1 0.71 1.035 0.71 1.035 0.675 0.895 0.675 0.895 0.905 0.86 0.905 0.86 1.045 0.795 1.045  ;
  END
END OAI21_X4

MACRO SDFFS_X1
  CLASS core ;
  FOREIGN SDFFS_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 5.51 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 4.98 0.42 5.08 0.42 5.08 0.985 4.98 0.985  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 3.02 0.4 3.085 0.4 3.085 0.435 3.23 0.435 3.23 0.175 3.465 0.175 3.465 0.16 3.565 0.16 3.565 0.175 4.295 0.175 4.295 0.545 4.44 0.545 4.44 0.51 4.505 0.51 4.505 0.645 4.44 0.645 4.44 0.61 4.23 0.61 4.23 0.24 3.565 0.24 3.565 0.26 3.465 0.26 3.465 0.24 3.295 0.24 3.295 0.5 3.085 0.5 3.085 0.535 3.02 0.535  ;
    END
  END SN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.425 0.62 0.525 0.62 0.525 0.755 0.425 0.755  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.335 1.315 0.335 1 0.4 1 0.4 1.315 1.095 1.315 1.095 1 1.16 1 1.16 1.315 1.655 1.315 1.655 1.025 1.72 1.025 1.72 1.315 2.09 1.315 2.09 1.025 2.155 1.025 2.155 1.315 2.865 1.315 2.865 1.125 2.93 1.125 2.93 1.315 3.42 1.315 3.42 1.09 3.485 1.09 3.485 1.315 4.36 1.315 4.36 1.05 4.425 1.05 4.425 1.315 4.735 1.315 4.735 1.015 4.8 1.015 4.8 1.315 5.165 1.315 5.165 0.91 5.23 0.91 5.23 1.315 5.51 1.315 5.51 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 5.32 0.42 5.42 0.42 5.42 0.985 5.32 0.985  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.385 0.49 0.425 0.49 0.425 0.44 0.525 0.44 0.525 0.49 0.96 0.49 0.96 0.455 1.025 0.455 1.025 0.59 0.96 0.59 0.96 0.555 0.385 0.555  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 5.51 -0.085 5.51 0.085 5.235 0.085 5.235 0.54 5.17 0.54 5.17 0.085 4.425 0.085 4.425 0.43 4.36 0.43 4.36 0.085 3.165 0.085 3.165 0.335 3.1 0.335 3.1 0.085 2.165 0.085 2.165 0.395 2.1 0.395 2.1 0.085 1.72 0.085 1.72 0.2 1.655 0.2 1.655 0.085 1.285 0.085 1.285 0.325 1.22 0.325 1.22 0.085 0.4 0.085 0.4 0.325 0.335 0.325 0.335 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.385 0.82 0.59 0.82 0.59 0.655 1.12 0.655 1.12 0.52 1.185 0.52 1.185 0.72 0.905 0.72 0.905 0.82 0.805 0.82 0.805 0.72 0.655 0.72 0.655 0.885 0.385 0.885  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.565 0.795 1.7 0.795 1.7 0.895 1.565 0.895  ;
    END
  END CK
  OBS
      LAYER M1 ;
        POLYGON 0.095 0.295 0.215 0.295 0.215 1.08 0.095 1.08  ;
        POLYGON 2.425 0.76 3.125 0.76 3.125 0.73 3.26 0.73 3.26 0.795 3.225 0.795 3.225 0.83 2.615 0.83 2.615 0.895 2.55 0.895 2.55 0.825 2.36 0.825 2.36 0.5 2.395 0.5 2.395 0.465 2.46 0.465 2.46 0.6 2.425 0.6  ;
        POLYGON 2.805 0.455 2.905 0.455 2.905 0.6 3.36 0.6 3.36 0.42 3.425 0.42 3.425 0.76 3.485 0.76 3.485 0.895 3.42 0.895 3.42 0.86 3.36 0.86 3.36 0.665 2.84 0.665 2.84 0.59 2.805 0.59  ;
        POLYGON 2.295 0.96 2.565 0.96 2.565 0.995 3.24 0.995 3.24 0.96 3.575 0.96 3.575 0.375 3.64 0.375 3.64 0.84 3.675 0.84 3.675 1.025 3.305 1.025 3.305 1.095 3.24 1.095 3.24 1.06 2.23 1.06 2.23 0.33 2.515 0.33 2.515 0.295 2.58 0.295 2.58 0.43 2.515 0.43 2.515 0.395 2.295 0.395  ;
        POLYGON 3.77 0.375 3.835 0.375 3.835 0.875 4.075 0.875 4.075 0.94 3.77 0.94  ;
        POLYGON 3.91 1.04 3.945 1.04 3.945 1.005 4.14 1.005 4.14 0.81 3.945 0.81 3.945 0.305 4.01 0.305 4.01 0.745 4.59 0.745 4.59 0.71 4.725 0.71 4.725 0.775 4.69 0.775 4.69 0.81 4.205 0.81 4.205 1.07 4.045 1.07 4.045 1.105 3.91 1.105  ;
        POLYGON 4.27 0.875 4.79 0.875 4.79 0.645 4.735 0.645 4.735 0.21 4.89 0.21 4.89 0.94 4.61 0.94 4.61 1.135 4.545 1.135 4.545 0.94 4.27 0.94  ;
        POLYGON 1.4 0.76 1.5 0.76 1.5 1.055 1.4 1.055  ;
        POLYGON 1.38 0.5 1.415 0.5 1.415 0.17 1.535 0.17 1.535 0.365 1.81 0.365 1.81 0.43 1.535 0.43 1.535 0.565 1.38 0.565  ;
        POLYGON 1.845 0.76 1.965 0.76 1.965 1.055 1.845 1.055  ;
        POLYGON 1.875 0.17 1.975 0.17 1.975 0.565 1.875 0.565  ;
        POLYGON 0.685 0.98 0.965 0.98 0.965 0.87 1.25 0.87 1.25 0.455 1.09 0.455 1.09 0.39 0.685 0.39 0.685 0.325 1.155 0.325 1.155 0.39 1.315 0.39 1.315 0.63 2.1 0.63 2.1 0.465 2.165 0.465 2.165 0.895 2.1 0.895 2.1 0.695 1.315 0.695 1.315 0.935 1.03 0.935 1.03 1.045 0.685 1.045  ;
  END
END SDFFS_X1

MACRO SDFFS_X2
  CLASS core ;
  FOREIGN SDFFS_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 5.51 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 4.98 0.42 5.08 0.42 5.08 0.985 4.98 0.985  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 3.02 0.4 3.085 0.4 3.085 0.435 3.23 0.435 3.23 0.175 3.465 0.175 3.465 0.16 3.565 0.16 3.565 0.175 4.295 0.175 4.295 0.545 4.44 0.545 4.44 0.51 4.505 0.51 4.505 0.645 4.44 0.645 4.44 0.61 4.23 0.61 4.23 0.24 3.565 0.24 3.565 0.26 3.465 0.26 3.465 0.24 3.295 0.24 3.295 0.5 3.085 0.5 3.085 0.535 3.02 0.535  ;
    END
  END SN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.425 0.62 0.525 0.62 0.525 0.755 0.425 0.755  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.335 1.315 0.335 1 0.4 1 0.4 1.315 1.095 1.315 1.095 1 1.16 1 1.16 1.315 1.655 1.315 1.655 1.025 1.72 1.025 1.72 1.315 2.09 1.315 2.09 1.025 2.155 1.025 2.155 1.315 2.865 1.315 2.865 1.125 2.93 1.125 2.93 1.315 3.42 1.315 3.42 1.09 3.485 1.09 3.485 1.315 4.36 1.315 4.36 1.05 4.425 1.05 4.425 1.315 4.735 1.315 4.735 1.015 4.8 1.015 4.8 1.315 5.165 1.315 5.165 1.045 5.23 1.045 5.23 1.315 5.51 1.315 5.51 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 5.32 0.42 5.42 0.42 5.42 0.985 5.32 0.985  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.385 0.49 0.425 0.49 0.425 0.44 0.525 0.44 0.525 0.49 0.96 0.49 0.96 0.455 1.025 0.455 1.025 0.59 0.96 0.59 0.96 0.555 0.385 0.555  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 5.51 -0.085 5.51 0.085 5.235 0.085 5.235 0.45 5.17 0.45 5.17 0.085 4.425 0.085 4.425 0.43 4.36 0.43 4.36 0.085 3.165 0.085 3.165 0.335 3.1 0.335 3.1 0.085 2.165 0.085 2.165 0.395 2.1 0.395 2.1 0.085 1.72 0.085 1.72 0.2 1.655 0.2 1.655 0.085 1.285 0.085 1.285 0.325 1.22 0.325 1.22 0.085 0.4 0.085 0.4 0.325 0.335 0.325 0.335 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.385 0.82 0.59 0.82 0.59 0.655 1.12 0.655 1.12 0.52 1.185 0.52 1.185 0.72 0.655 0.72 0.655 0.885 0.385 0.885  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.565 0.795 1.7 0.795 1.7 0.895 1.565 0.895  ;
    END
  END CK
  OBS
      LAYER M1 ;
        POLYGON 0.095 0.295 0.215 0.295 0.215 1.08 0.095 1.08  ;
        POLYGON 2.425 0.76 3.125 0.76 3.125 0.73 3.26 0.73 3.26 0.795 3.225 0.795 3.225 0.83 2.615 0.83 2.615 0.895 2.55 0.895 2.55 0.825 2.36 0.825 2.36 0.5 2.395 0.5 2.395 0.465 2.46 0.465 2.46 0.6 2.425 0.6  ;
        POLYGON 2.805 0.455 2.905 0.455 2.905 0.6 3.36 0.6 3.36 0.42 3.425 0.42 3.425 0.76 3.485 0.76 3.485 0.895 3.42 0.895 3.42 0.86 3.36 0.86 3.36 0.665 2.84 0.665 2.84 0.59 2.805 0.59  ;
        POLYGON 2.295 0.96 2.565 0.96 2.565 0.995 3.24 0.995 3.24 0.96 3.575 0.96 3.575 0.375 3.64 0.375 3.64 0.84 3.675 0.84 3.675 1.025 3.305 1.025 3.305 1.095 3.24 1.095 3.24 1.06 2.23 1.06 2.23 0.33 2.515 0.33 2.515 0.295 2.58 0.295 2.58 0.43 2.515 0.43 2.515 0.395 2.295 0.395  ;
        POLYGON 3.77 0.375 3.835 0.375 3.835 0.87 4.075 0.87 4.075 0.935 3.77 0.935  ;
        POLYGON 3.91 1.035 3.945 1.035 3.945 1 4.14 1 4.14 0.78 3.945 0.78 3.945 0.305 4.01 0.305 4.01 0.715 4.565 0.715 4.565 0.68 4.7 0.68 4.7 0.745 4.665 0.745 4.665 0.78 4.205 0.78 4.205 1.065 4.045 1.065 4.045 1.1 3.91 1.1  ;
        POLYGON 4.27 0.875 4.79 0.875 4.79 0.645 4.755 0.645 4.755 0.21 4.89 0.21 4.89 0.94 4.615 0.94 4.615 1.135 4.55 1.135 4.55 0.94 4.27 0.94  ;
        POLYGON 1.4 0.76 1.5 0.76 1.5 1.055 1.4 1.055  ;
        POLYGON 1.38 0.5 1.415 0.5 1.415 0.17 1.535 0.17 1.535 0.365 1.81 0.365 1.81 0.43 1.535 0.43 1.535 0.565 1.38 0.565  ;
        POLYGON 1.845 0.76 1.965 0.76 1.965 1.055 1.845 1.055  ;
        POLYGON 1.875 0.17 1.975 0.17 1.975 0.565 1.875 0.565  ;
        POLYGON 0.685 0.98 0.755 0.98 0.755 0.87 1.25 0.87 1.25 0.455 1.09 0.455 1.09 0.39 0.685 0.39 0.685 0.325 1.155 0.325 1.155 0.39 1.315 0.39 1.315 0.63 2.1 0.63 2.1 0.465 2.165 0.465 2.165 0.895 2.1 0.895 2.1 0.695 1.315 0.695 1.315 0.935 0.82 0.935 0.82 1.045 0.685 1.045  ;
  END
END SDFFS_X2

MACRO SDFFR_X1
  CLASS core ;
  FOREIGN SDFFR_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 5.51 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.42 0.185 0.42 0.185 1.03 0.05 1.03  ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 4.795 0.62 4.895 0.62 4.895 0.755 4.795 0.755  ;
    END
  END SE
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.49 0.86 1.625 0.86 1.625 0.895 1.755 0.895 1.755 0.86 1.855 0.86 1.855 0.895 2.055 0.895 2.055 0.86 2.825 0.86 2.825 0.995 2.76 0.995 2.76 0.925 2.115 0.925 2.115 0.96 1.855 0.96 1.755 0.96 1.525 0.96 1.525 0.925 1.49 0.925  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.27 1.315 0.27 1.02 0.27 0.955 0.335 0.955 0.335 1.315 0.875 1.315 0.875 1.08 0.94 1.08 0.94 1.315 1.635 1.315 1.635 1.17 1.7 1.17 1.7 1.315 2.515 1.315 2.515 1.06 2.58 1.06 2.58 1.315 3.02 1.315 3.02 1.1 3.085 1.1 3.085 1.315 3.81 1.315 3.81 1.1 3.875 1.1 3.875 1.315 4.325 1.315 4.325 1 4.39 1 4.39 1.315 5.08 1.315 5.08 1 5.145 1 5.145 1.315 5.51 1.315 5.51 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.425 0.42 0.56 0.42 0.56 1.03 0.425 1.03  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 4.425 0.61 4.46 0.61 4.46 0.49 5 0.49 5 0.455 5.065 0.455 5.065 0.59 5 0.59 5 0.555 4.56 0.555 4.56 0.675 4.425 0.675  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 5.51 -0.085 5.51 0.085 5.15 0.085 5.15 0.15 5.15 0.325 5.085 0.325 5.085 0.085 4.275 0.085 4.275 0.325 4.21 0.325 4.21 0.085 3.875 0.085 3.875 0.265 3.81 0.265 3.81 0.085 3.08 0.085 3.08 0.265 3.015 0.265 3.015 0.085 1.89 0.085 1.89 0.36 1.825 0.36 1.825 0.085 0.94 0.085 0.94 0.36 0.875 0.36 0.875 0.085 0.335 0.085 0.335 0.54 0.27 0.54 0.27 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 4.295 0.52 4.36 0.52 4.36 0.74 4.65 0.74 4.65 0.82 5 0.82 5 0.785 5.065 0.785 5.065 0.92 5 0.92 5 0.885 4.585 0.885 4.585 0.805 4.295 0.805  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 3.885 0.705 3.985 0.705 3.985 0.84 3.885 0.84  ;
    END
  END CK
  OBS
      LAYER M1 ;
        POLYGON 3.665 0.905 4.1 0.905 4.1 1.04 4 1.04 4 0.97 3.665 0.97 3.665 1.225 3.27 1.225 3.27 0.865 3.235 0.865 3.235 0.83 2.885 0.83 2.885 0.795 1.995 0.795 1.995 0.83 1.93 0.83 1.93 0.685 1.505 0.685 1.505 0.72 1.44 0.72 1.44 0.585 1.505 0.585 1.505 0.62 1.995 0.62 1.995 0.73 2.365 0.73 2.365 0.62 2.5 0.62 2.5 0.73 2.945 0.73 2.945 0.765 3.235 0.765 3.235 0.73 3.3 0.73 3.3 0.765 3.335 0.765 3.335 1.16 3.6 1.16 3.6 0.53 3.565 0.53 3.565 0.395 3.6 0.395 3.6 0.33 3.965 0.33 3.965 0.235 4.065 0.235 4.065 0.395 3.665 0.395  ;
        POLYGON 3.73 0.46 3.795 0.46 3.795 0.495 4.165 0.495 4.165 0.39 4.34 0.39 4.34 0.33 4.8 0.33 4.8 0.395 4.405 0.395 4.405 0.455 4.23 0.455 4.23 0.87 4.52 0.87 4.52 0.95 4.765 0.95 4.765 1.085 4.7 1.085 4.7 1.015 4.455 1.015 4.455 0.935 4.165 0.935 4.165 0.56 3.795 0.56 3.795 0.595 3.73 0.595  ;
        POLYGON 5.27 0.295 5.39 0.295 5.39 1.08 5.27 1.08  ;
        POLYGON 0.65 0.28 0.75 0.28 0.75 1.2 0.65 1.2  ;
        POLYGON 1.245 1.08 1.315 1.08 1.315 1.15 1.505 1.15 1.505 1.04 1.83 1.04 1.83 1.115 2.01 1.115 2.01 1.08 2.075 1.08 2.075 1.215 2.01 1.215 2.01 1.18 1.765 1.18 1.765 1.105 1.57 1.105 1.57 1.215 1.25 1.215 1.25 1.18 1.18 1.18 1.18 0.715 0.88 0.715 0.88 1.015 0.815 1.015 0.815 0.58 0.88 0.58 0.88 0.65 1.18 0.65 1.18 0.27 1.54 0.27 1.54 0.335 1.245 0.335  ;
        POLYGON 2.17 0.995 2.235 0.995 2.235 1.03 2.33 1.03 2.33 0.995 2.395 0.995 2.395 1.13 2.33 1.13 2.33 1.095 2.235 1.095 2.235 1.13 2.17 1.13  ;
        POLYGON 2.605 0.18 2.95 0.18 2.95 0.34 3.2 0.34 3.2 0.405 2.885 0.405 2.885 0.245 2.605 0.245  ;
        POLYGON 2.83 1.06 2.89 1.06 2.89 0.96 3.14 0.96 3.14 0.925 3.205 0.925 3.205 1.06 3.14 1.06 3.14 1.025 2.955 1.025 2.955 1.16 2.895 1.16 2.895 1.195 2.83 1.195  ;
        POLYGON 1.31 0.4 1.615 0.4 1.615 0.47 2.01 0.47 2.01 0.33 2.075 0.33 2.075 0.365 2.235 0.365 2.235 0.435 2.82 0.435 2.82 0.47 3.305 0.47 3.305 0.4 3.37 0.4 3.37 0.535 2.76 0.535 2.76 0.5 2.07 0.5 2.07 0.535 1.55 0.535 1.55 0.5 1.375 0.5 1.375 1.015 1.31 1.015  ;
        POLYGON 3.4 1.03 3.47 1.03 3.47 0.665 2.6 0.665 2.6 0.63 2.565 0.63 2.565 0.565 2.7 0.565 2.7 0.6 3.435 0.6 3.435 0.15 3.5 0.15 3.5 0.605 3.535 0.605 3.535 1.095 3.4 1.095  ;
  END
END SDFFR_X1

MACRO SDFFR_X2
  CLASS core ;
  FOREIGN SDFFR_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 5.51 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.42 0.15 0.42 0.15 1.17 0.05 1.17  ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 4.795 0.62 4.895 0.62 4.895 0.755 4.795 0.755  ;
    END
  END SE
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.49 0.86 1.625 0.86 1.625 0.895 1.755 0.895 1.755 0.86 1.855 0.86 1.855 0.895 2.055 0.895 2.055 0.86 2.825 0.86 2.825 0.995 2.76 0.995 2.76 0.925 2.115 0.925 2.115 0.96 1.855 0.96 1.755 0.96 1.525 0.96 1.525 0.925 1.49 0.925  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.27 1.315 0.27 1.015 0.27 0.95 0.335 0.95 0.335 1.315 0.875 1.315 0.875 1.095 0.94 1.095 0.94 1.315 1.635 1.315 1.635 1.185 1.7 1.185 1.7 1.315 2.515 1.315 2.515 1.06 2.58 1.06 2.58 1.315 3.02 1.315 3.02 1.1 3.085 1.1 3.085 1.315 3.81 1.315 3.81 1.1 3.875 1.1 3.875 1.315 4.315 1.315 4.315 1 4.38 1 4.38 1.315 5.07 1.315 5.07 1 5.135 1 5.135 1.315 5.51 1.315 5.51 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.425 0.42 0.56 0.42 0.56 1.17 0.425 1.17  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 4.415 0.61 4.45 0.61 4.45 0.49 4.99 0.49 4.99 0.455 5.055 0.455 5.055 0.59 4.99 0.59 4.99 0.555 4.55 0.555 4.55 0.675 4.415 0.675  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 5.51 -0.085 5.51 0.085 5.14 0.085 5.14 0.15 5.14 0.325 5.075 0.325 5.075 0.085 4.265 0.085 4.265 0.325 4.2 0.325 4.2 0.085 3.875 0.085 3.875 0.265 3.81 0.265 3.81 0.085 3.08 0.085 3.08 0.265 3.015 0.265 3.015 0.085 1.89 0.085 1.89 0.36 1.825 0.36 1.825 0.085 0.94 0.085 0.94 0.36 0.875 0.36 0.875 0.085 0.335 0.085 0.335 0.45 0.27 0.45 0.27 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 4.285 0.52 4.35 0.52 4.35 0.74 4.64 0.74 4.64 0.82 4.99 0.82 4.99 0.785 5.055 0.785 5.055 0.92 4.99 0.92 4.99 0.885 4.575 0.885 4.575 0.805 4.285 0.805  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 3.885 0.685 3.985 0.685 3.985 0.82 3.885 0.82  ;
    END
  END CK
  OBS
      LAYER M1 ;
        POLYGON 3.665 0.97 4.1 0.97 4.1 1.105 4 1.105 4 1.035 3.665 1.035 3.665 1.225 3.27 1.225 3.27 0.865 3.235 0.865 3.235 0.83 2.885 0.83 2.885 0.795 1.995 0.795 1.995 0.83 1.93 0.83 1.93 0.7 1.53 0.7 1.53 0.735 1.465 0.735 1.465 0.6 1.53 0.6 1.53 0.635 1.995 0.635 1.995 0.73 2.365 0.73 2.365 0.635 2.5 0.635 2.5 0.73 2.945 0.73 2.945 0.765 3.235 0.765 3.235 0.73 3.3 0.73 3.3 0.765 3.335 0.765 3.335 1.16 3.6 1.16 3.6 0.53 3.565 0.53 3.565 0.395 3.6 0.395 3.6 0.33 3.965 0.33 3.965 0.235 4.065 0.235 4.065 0.395 3.665 0.395  ;
        POLYGON 3.73 0.46 3.795 0.46 3.795 0.495 4.155 0.495 4.155 0.39 4.33 0.39 4.33 0.33 4.79 0.33 4.79 0.395 4.395 0.395 4.395 0.455 4.22 0.455 4.22 0.87 4.51 0.87 4.51 0.95 4.755 0.95 4.755 1.085 4.69 1.085 4.69 1.015 4.445 1.015 4.445 0.935 4.155 0.935 4.155 0.56 3.795 0.56 3.795 0.595 3.73 0.595  ;
        POLYGON 5.26 0.295 5.38 0.295 5.38 1.08 5.26 1.08  ;
        POLYGON 0.65 0.28 0.75 0.28 0.75 1.215 0.65 1.215  ;
        POLYGON 1.27 1.095 1.315 1.095 1.315 1.165 1.505 1.165 1.505 1.055 1.83 1.055 1.83 1.13 2.01 1.13 2.01 1.095 2.075 1.095 2.075 1.23 2.01 1.23 2.01 1.195 1.765 1.195 1.765 1.12 1.57 1.12 1.57 1.23 1.25 1.23 1.25 1.195 1.205 1.195 1.205 0.715 0.88 0.715 0.88 1.03 0.815 1.03 0.815 0.58 0.88 0.58 0.88 0.65 1.205 0.65 1.205 0.27 1.54 0.27 1.54 0.335 1.27 0.335  ;
        POLYGON 2.17 0.995 2.235 0.995 2.235 1.03 2.33 1.03 2.33 0.995 2.395 0.995 2.395 1.13 2.33 1.13 2.33 1.095 2.235 1.095 2.235 1.13 2.17 1.13  ;
        POLYGON 2.605 0.18 2.95 0.18 2.95 0.34 3.2 0.34 3.2 0.405 2.885 0.405 2.885 0.245 2.605 0.245  ;
        POLYGON 2.83 1.06 2.89 1.06 2.89 0.96 3.14 0.96 3.14 0.925 3.205 0.925 3.205 1.06 3.14 1.06 3.14 1.025 2.955 1.025 2.955 1.16 2.895 1.16 2.895 1.195 2.83 1.195  ;
        POLYGON 1.335 0.4 1.615 0.4 1.615 0.465 2.01 0.465 2.01 0.33 2.075 0.33 2.075 0.365 2.235 0.365 2.235 0.435 2.82 0.435 2.82 0.47 3.305 0.47 3.305 0.4 3.37 0.4 3.37 0.535 2.76 0.535 2.76 0.5 2.065 0.5 2.065 0.535 1.4 0.535 1.4 1.03 1.335 1.03  ;
        POLYGON 3.4 1.03 3.47 1.03 3.47 0.665 2.6 0.665 2.6 0.63 2.565 0.63 2.565 0.565 2.7 0.565 2.7 0.6 3.435 0.6 3.435 0.15 3.5 0.15 3.5 0.605 3.535 0.605 3.535 1.095 3.4 1.095  ;
  END
END SDFFR_X2

MACRO DFFSRX1  #DFFRS_X1
  CLASS core ;
  #FOREIGN DFFRS_X1 0.0 0.0 ;
  FOREIGN DFFSRX1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 5.89 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 5.755 0.735 5.79 0.735 5.79 0.4 5.745 0.4 5.745 0.3 5.755 0.3 5.755 0.285 5.755 0.15 5.82 0.15 5.82 0.185 5.855 0.185 5.855 0.835 5.82 0.835 5.82 0.87 5.755 0.87  ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
	CAPACITANCE 0.007439 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 4.01 0.75 4.455 0.75 4.455 0.955 4.39 0.955 4.39 0.815 3.945 0.815 3.945 0.65 3.91 0.65 3.91 0.585 3.945 0.585 3.945 0.425 3.645 0.425 3.645 0.27 2.885 0.27 2.885 0.425 2.49 0.425 2.49 0.27 2.095 0.27 2.095 0.59 1.75 0.59 1.75 0.525 2.03 0.525 2.03 0.205 2.135 0.205 2.135 0.16 2.235 0.16 2.235 0.205 2.555 0.205 2.555 0.36 2.82 0.36 2.82 0.205 3.71 0.205 3.71 0.36 4.01 0.36 4.01 0.585 4.045 0.585 4.045 0.65 4.01 0.65  ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
	CAPACITANCE 0.001967 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 2.8 0.755 3.075 0.755 3.075 0.72 3.275 0.72 3.375 0.72 3.715 0.72 3.715 0.785 3.375 0.785 3.375 0.82 3.275 0.82 3.275 0.785 3.135 0.785 3.135 0.82 2.8 0.82  ;
    END
  END SN
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 3.42 1.315 4.13 1.315 4.13 1.06 4.195 1.06 4.195 1.315 4.85 1.315 4.85 0.685 4.95 0.685 4.95 1.315 5.23 1.315 5.23 0.685 5.295 0.685 5.295 1.315 5.57 1.315 5.57 0.795 5.635 0.795 5.635 1.315 5.89 1.315 5.89 1.485 0 1.485 0 1.315 0.275 1.315 0.275 0.9 0.34 0.9 0.34 1.315 1.03 1.315 1.03 1.155 1.095 1.155 1.095 1.315 1.89 1.315 1.89 1.075 1.955 1.075 1.955 1.315 2.635 1.315 2.635 1.13 2.6 1.13 2.6 1.065 2.735 1.065 2.735 1.13 2.7 1.13 2.7 1.315 3.355 1.315 3.355 1.175 3.32 1.175 3.32 1.11 3.455 1.11 3.455 1.175 3.42 1.175  ;
    END
  END POWR  #VDD
  PIN Q
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 5.365 0.72 5.415 0.72 5.415 0.665 5.6 0.665 5.6 0.4 5.415 0.4 5.415 0.265 5.48 0.265 5.48 0.335 5.665 0.335 5.665 0.73 5.48 0.73 5.48 0.8 5.465 0.8 5.465 0.82 5.365 0.82  ;
    END
  END Q
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 3.775 0.23 3.81 0.23 3.81 0.085 2.72 0.085 2.72 0.23 2.755 0.23 2.755 0.295 2.62 0.295 2.62 0.23 2.655 0.23 2.655 0.085 1.93 0.085 1.93 0.35 1.965 0.35 1.965 0.415 1.83 0.415 1.83 0.35 1.865 0.35 1.865 0.085 0.7 0.085 0.7 0.36 0.635 0.36 0.635 0.085 0.34 0.085 0.34 0.355 0.275 0.355 0.275 0.15 0.275 0.085 0 0.085 0 -0.085 5.89 -0.085 5.89 0.085 5.635 0.085 5.635 0.27 5.57 0.27 5.57 0.085 5.295 0.085 5.295 0.4 5.23 0.4 5.23 0.085 3.875 0.085 3.875 0.23 3.91 0.23 3.91 0.295 3.775 0.295  ;
    END
  END GRND  #VSS
  PIN D
    DIRECTION INPUT ;
	CAPACITANCE 0.000958 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.615 0.545 0.715 0.545 0.715 0.68 0.615 0.68  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
	CAPACITANCE 0.000515 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.205 0.685 0.34 0.685 0.34 0.82 0.205 0.82  ;
    END
  END CK
  OBS
      LAYER M1 ;
        POLYGON 0.04 0.325 0.155 0.325 0.155 0.52 0.35 0.52 0.35 0.485 0.415 0.485 0.415 0.62 0.35 0.62 0.35 0.585 0.14 0.585 0.14 1.12 0.04 1.12  ;
        POLYGON 2.735 0.935 2.955 0.935 2.955 0.97 3.585 0.97 3.585 1.04 4 1.04 4 0.93 4.325 0.93 4.325 1.02 4.555 1.02 4.555 0.945 4.52 0.945 4.52 0.88 4.555 0.88 4.555 0.685 4.11 0.685 4.11 0.55 4.175 0.55 4.175 0.62 4.62 0.62 4.62 0.88 4.655 0.88 4.655 0.945 4.62 0.945 4.62 1.085 4.26 1.085 4.26 0.995 4.065 0.995 4.065 1.105 3.52 1.105 3.52 1.035 2.855 1.035 2.855 1 2.67 1 2.67 0.625 2.95 0.625 2.95 0.335 3.165 0.335 3.165 0.4 3.015 0.4 3.015 0.69 2.735 0.69  ;
        POLYGON 4.415 1.15 4.72 1.15 4.72 0.295 4.41 0.295 4.41 0.33 4.345 0.33 4.345 0.295 4.15 0.295 4.15 0.23 4.345 0.23 4.345 0.195 4.41 0.195 4.41 0.23 4.785 0.23 4.785 1.215 4.415 1.215  ;
        POLYGON 4.85 0.32 4.915 0.32 4.915 0.5 5.47 0.5 5.47 0.465 5.535 0.465 5.535 0.6 5.47 0.6 5.47 0.565 5.1 0.565 5.1 0.76 5.035 0.76 5.035 0.565 4.85 0.565  ;
        POLYGON 0.48 0.325 0.545 0.325 0.545 0.745 0.95 0.745 0.95 0.71 1.015 0.71 1.015 0.845 0.95 0.845 0.95 0.81 0.545 0.81 0.545 0.98 0.48 0.98  ;
        POLYGON 1.28 0.81 1.315 0.81 1.315 0.595 0.86 0.595 0.86 0.53 1.38 0.53 1.38 0.81 1.415 0.81 1.415 0.875 1.28 0.875  ;
        POLYGON 0.655 0.875 0.72 0.875 0.72 1.005 1.48 1.005 1.48 0.43 1.365 0.43 1.365 0.465 1.3 0.465 1.3 0.33 1.365 0.33 1.365 0.365 1.545 0.365 1.545 0.935 2.35 0.935 2.35 1.145 2.285 1.145 2.285 1 1.58 1 1.58 1.21 1.515 1.21 1.515 1.07 0.72 1.07 0.72 1.15 0.655 1.15  ;
        POLYGON 1.61 0.655 2.23 0.655 2.23 0.4 2.16 0.4 2.16 0.335 2.295 0.335 2.295 0.665 2.48 0.665 2.48 0.835 2.515 0.835 2.515 1.11 2.45 1.11 2.45 0.97 2.415 0.97 2.415 0.73 2.26 0.73 2.26 0.72 1.61 0.72  ;
        POLYGON 2.36 0.495 2.885 0.495 2.885 0.56 2.36 0.56  ;
        POLYGON 3.08 0.495 3.215 0.495 3.215 0.535 3.845 0.535 3.845 0.88 3.915 0.88 3.915 0.945 3.78 0.945 3.78 0.6 3.155 0.6 3.155 0.56 3.08 0.56  ;
  END
END DFFSRX1  #DFFRS_X1

MACRO DFFRS_X2
  CLASS core ;
  FOREIGN DFFRS_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 6.08 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 5.77 0.74 5.805 0.74 5.805 0.54 5.745 0.54 5.745 0.44 5.805 0.44 5.805 0.375 5.77 0.375 5.77 0.24 5.835 0.24 5.835 0.275 5.87 0.275 5.87 0.875 5.835 0.875 5.835 1.015 5.77 1.015  ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 4.01 0.75 4.455 0.75 4.455 0.955 4.39 0.955 4.39 0.815 3.945 0.815 3.945 0.65 3.91 0.65 3.91 0.585 3.945 0.585 3.945 0.425 3.645 0.425 3.645 0.27 2.885 0.27 2.885 0.425 2.49 0.425 2.49 0.27 2.095 0.27 2.095 0.59 1.75 0.59 1.75 0.525 2.03 0.525 2.03 0.205 2.135 0.205 2.135 0.16 2.235 0.16 2.235 0.205 2.555 0.205 2.555 0.36 2.82 0.36 2.82 0.205 3.71 0.205 3.71 0.36 4.01 0.36 4.01 0.585 4.045 0.585 4.045 0.65 4.01 0.65  ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 2.8 0.755 3.075 0.755 3.075 0.72 3.275 0.72 3.375 0.72 3.715 0.72 3.715 0.785 3.375 0.785 3.375 0.82 3.275 0.82 3.275 0.785 3.135 0.785 3.135 0.82 2.8 0.82  ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 3.42 1.315 4.13 1.315 4.13 1.06 4.195 1.06 4.195 1.315 4.85 1.315 4.85 0.685 4.95 0.685 4.95 1.315 5.245 1.315 5.245 0.68 5.31 0.68 5.31 1.315 5.585 1.315 5.585 0.795 5.65 0.795 5.65 1.315 6.08 1.315 6.08 1.485 0 1.485 0 1.315 0.275 1.315 0.275 0.9 0.34 0.9 0.34 1.315 1.03 1.315 1.03 1.155 1.095 1.155 1.095 1.315 1.89 1.315 1.89 1.075 1.955 1.075 1.955 1.315 2.635 1.315 2.635 1.13 2.6 1.13 2.6 1.065 2.735 1.065 2.735 1.13 2.7 1.13 2.7 1.315 3.355 1.315 3.355 1.175 3.32 1.175 3.32 1.11 3.455 1.11 3.455 1.175 3.42 1.175  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 5.43 0.665 5.615 0.665 5.615 0.4 5.43 0.4 5.43 0.265 5.495 0.265 5.495 0.335 5.68 0.335 5.68 0.73 5.495 0.73 5.495 0.94 5.43 0.94  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 3.775 0.23 3.81 0.23 3.81 0.085 2.72 0.085 2.72 0.23 2.755 0.23 2.755 0.295 2.62 0.295 2.62 0.23 2.655 0.23 2.655 0.085 1.93 0.085 1.93 0.35 1.965 0.35 1.965 0.415 1.83 0.415 1.83 0.35 1.865 0.35 1.865 0.085 0.7 0.085 0.7 0.36 0.635 0.36 0.635 0.085 0.34 0.085 0.34 0.355 0.275 0.355 0.275 0.15 0.275 0.085 0 0.085 0 -0.085 6.08 -0.085 6.08 0.085 5.65 0.085 5.65 0.27 5.585 0.27 5.585 0.085 5.31 0.085 5.31 0.335 5.245 0.335 5.245 0.085 3.875 0.085 3.875 0.23 3.91 0.23 3.91 0.295 3.775 0.295  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.615 0.545 0.715 0.545 0.715 0.68 0.615 0.68  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.205 0.685 0.34 0.685 0.34 0.82 0.205 0.82  ;
    END
  END CK
  OBS
      LAYER M1 ;
        POLYGON 0.04 0.325 0.155 0.325 0.155 0.52 0.35 0.52 0.35 0.485 0.415 0.485 0.415 0.62 0.35 0.62 0.35 0.585 0.14 0.585 0.14 1.12 0.04 1.12  ;
        POLYGON 2.735 0.935 2.955 0.935 2.955 0.97 3.585 0.97 3.585 1.04 4 1.04 4 0.93 4.325 0.93 4.325 1.02 4.555 1.02 4.555 0.945 4.52 0.945 4.52 0.88 4.555 0.88 4.555 0.685 4.11 0.685 4.11 0.55 4.175 0.55 4.175 0.62 4.62 0.62 4.62 0.88 4.655 0.88 4.655 0.945 4.62 0.945 4.62 1.085 4.26 1.085 4.26 0.995 4.065 0.995 4.065 1.105 3.52 1.105 3.52 1.035 2.855 1.035 2.855 1 2.67 1 2.67 0.625 2.95 0.625 2.95 0.335 3.165 0.335 3.165 0.4 3.015 0.4 3.015 0.69 2.735 0.69  ;
        POLYGON 4.415 1.15 4.72 1.15 4.72 0.295 4.41 0.295 4.41 0.33 4.345 0.33 4.345 0.295 4.15 0.295 4.15 0.23 4.345 0.23 4.345 0.195 4.41 0.195 4.41 0.23 4.785 0.23 4.785 1.215 4.415 1.215  ;
        POLYGON 4.85 0.305 4.915 0.305 4.915 0.5 5.485 0.5 5.485 0.465 5.55 0.465 5.55 0.6 5.485 0.6 5.485 0.565 5.1 0.565 5.1 0.76 5.035 0.76 5.035 0.565 4.85 0.565  ;
        POLYGON 0.48 0.325 0.545 0.325 0.545 0.745 0.95 0.745 0.95 0.71 1.015 0.71 1.015 0.845 0.95 0.845 0.95 0.81 0.545 0.81 0.545 0.98 0.48 0.98  ;
        POLYGON 1.28 0.81 1.315 0.81 1.315 0.595 0.86 0.595 0.86 0.53 1.38 0.53 1.38 0.81 1.415 0.81 1.415 0.875 1.28 0.875  ;
        POLYGON 0.655 0.875 0.72 0.875 0.72 1.005 1.48 1.005 1.48 0.43 1.365 0.43 1.365 0.465 1.3 0.465 1.3 0.33 1.365 0.33 1.365 0.365 1.545 0.365 1.545 0.935 2.35 0.935 2.35 1.145 2.285 1.145 2.285 1 1.58 1 1.58 1.21 1.515 1.21 1.515 1.07 0.72 1.07 0.72 1.15 0.655 1.15  ;
        POLYGON 1.61 0.655 2.23 0.655 2.23 0.4 2.16 0.4 2.16 0.335 2.295 0.335 2.295 0.665 2.48 0.665 2.48 0.835 2.515 0.835 2.515 1.11 2.45 1.11 2.45 0.97 2.415 0.97 2.415 0.73 2.26 0.73 2.26 0.72 1.61 0.72  ;
        POLYGON 2.36 0.495 2.885 0.495 2.885 0.56 2.36 0.56  ;
        POLYGON 3.08 0.495 3.215 0.495 3.215 0.535 3.845 0.535 3.845 0.88 3.915 0.88 3.915 0.945 3.78 0.945 3.78 0.6 3.155 0.6 3.155 0.56 3.08 0.56  ;
  END
END DFFRS_X2

MACRO DFFS_X1
  CLASS core ;
  FOREIGN DFFS_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 4.56 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 4.32 0.42 4.42 0.42 4.42 1.205 4.32 1.205  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.635 0.615 1.755 0.615 1.755 0.58 1.855 0.58 1.855 0.615 2.03 0.615 2.03 0.715 2.52 0.715 2.52 0.645 2.585 0.645 2.585 0.78 1.965 0.78 1.965 0.68 1.855 0.68 1.755 0.68 1.635 0.68  ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 3.4 1.315 4.13 1.315 4.13 1.13 4.195 1.13 4.195 1.315 4.56 1.315 4.56 1.485 0 1.485 0 1.315 0.235 1.315 0.235 0.82 0.3 0.82 0.3 1.315 0.61 1.315 0.61 0.995 0.675 0.995 0.675 1.315 1.48 1.315 1.48 1.07 1.545 1.07 1.545 1.315 1.91 1.315 1.91 0.985 1.975 0.985 1.975 1.315 2.485 1.315 2.485 1.17 2.45 1.17 2.45 1.105 2.585 1.105 2.585 1.17 2.55 1.17 2.55 1.315 3.335 1.315 3.335 1.17 3.3 1.17 3.3 1.105 3.435 1.105 3.435 1.17 3.4 1.17  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 3.89 0.42 4.01 0.42 4.01 0.715 3.89 0.715  ;
        POLYGON 3.89 0.91 4.01 0.91 4.01 1.205 3.89 1.205  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 2.375 0.255 2.41 0.255 2.41 0.085 1.445 0.085 1.445 0.445 1.38 0.445 1.38 0.085 0.675 0.085 0.675 0.355 0.61 0.355 0.61 0.085 0.3 0.085 0.3 0.275 0.235 0.275 0.235 0.085 0 0.085 0 -0.085 4.56 -0.085 4.56 0.085 4.195 0.085 4.195 0.54 4.13 0.54 4.13 0.085 3.59 0.085 3.59 0.39 3.525 0.39 3.525 0.085 2.475 0.085 2.475 0.255 2.51 0.255 2.51 0.32 2.375 0.32  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.615 0.615 0.715 0.615 0.715 0.75 0.615 0.75  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.18 0.605 0.315 0.605 0.315 0.74 0.18 0.74  ;
    END
  END CK
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.245 0.115 0.245 0.115 0.28 0.15 0.28 0.15 0.44 0.325 0.44 0.325 0.405 0.39 0.405 0.39 0.54 0.325 0.54 0.325 0.505 0.115 0.505 0.115 1.04 0.05 1.04  ;
        POLYGON 2.925 1.09 2.995 1.09 2.995 0.975 3.695 0.975 3.695 0.52 3.125 0.52 3.125 0.37 2.64 0.37 2.64 0.45 2.42 0.45 2.42 0.585 2.455 0.585 2.455 0.65 2.32 0.65 2.32 0.585 2.355 0.585 2.355 0.385 2.575 0.385 2.575 0.305 3.19 0.305 3.19 0.455 3.76 0.455 3.76 0.78 4.19 0.78 4.19 0.745 4.255 0.745 4.255 0.88 4.19 0.88 4.19 0.845 3.795 0.845 3.795 1.16 3.73 1.16 3.73 1.04 3.06 1.04 3.06 1.155 2.925 1.155  ;
        POLYGON 0.455 0.245 0.52 0.245 0.52 0.815 0.86 0.815 0.86 0.52 1.04 0.52 1.04 0.485 1.105 0.485 1.105 0.62 1.04 0.62 1.04 0.585 0.925 0.585 0.925 0.915 0.86 0.915 0.86 0.88 0.52 0.88 0.52 0.95 0.455 0.95  ;
        POLYGON 1.3 0.875 1.435 0.875 1.435 0.91 1.665 0.91 1.665 0.875 1.73 0.875 1.73 1.01 1.665 1.01 1.665 0.975 1.335 0.975 1.335 0.94 1.3 0.94  ;
        POLYGON 1.3 0.52 1.51 0.52 1.51 0.36 1.91 0.36 1.91 0.325 1.975 0.325 1.975 0.46 1.91 0.46 1.91 0.425 1.575 0.425 1.575 0.585 1.3 0.585  ;
        POLYGON 2.065 0.39 2.225 0.39 2.225 0.25 2.29 0.25 2.29 0.525 2.13 0.525 2.13 0.56 2.065 0.56  ;
        POLYGON 2.055 0.975 2.815 0.975 2.815 0.895 2.78 0.895 2.78 0.83 3.315 0.83 3.315 0.895 2.88 0.895 2.88 1.04 2.345 1.04 2.345 1.11 2.28 1.11 2.28 1.075 2.055 1.075  ;
        POLYGON 0.985 0.94 1.05 0.94 1.05 1.01 1.17 1.01 1.17 0.385 1.05 0.385 1.05 0.42 0.985 0.42 0.985 0.285 1.05 0.285 1.05 0.32 1.235 0.32 1.235 0.745 1.895 0.745 1.895 0.845 2.65 0.845 2.65 0.7 3.52 0.7 3.52 0.765 2.715 0.765 2.715 0.91 1.795 0.91 1.795 0.81 1.235 0.81 1.235 1.075 1.05 1.075 1.05 1.215 0.985 1.215  ;
  END
END DFFS_X1

MACRO DFFS_X2
  CLASS core ;
  FOREIGN DFFS_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 4.56 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 4.32 0.31 4.42 0.31 4.42 1.235 4.32 1.235  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.635 0.62 1.755 0.62 1.755 0.58 1.855 0.58 1.855 0.62 2.03 0.62 2.03 0.72 2.52 0.72 2.52 0.65 2.585 0.65 2.585 0.785 1.965 0.785 1.965 0.685 1.635 0.685  ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 3.405 1.315 4.13 1.315 4.13 1.015 4.195 1.015 4.195 1.315 4.56 1.315 4.56 1.485 0 1.485 0 1.315 0.235 1.315 0.235 0.825 0.3 0.825 0.3 1.315 0.61 1.315 0.61 1 0.675 1 0.675 1.315 1.48 1.315 1.48 1.075 1.545 1.075 1.545 1.315 1.91 1.315 1.91 0.99 1.975 0.99 1.975 1.315 2.485 1.315 2.485 1.175 2.45 1.175 2.45 1.11 2.585 1.11 2.585 1.175 2.55 1.175 2.55 1.315 3.34 1.315 3.34 1.175 3.305 1.175 3.305 1.11 3.44 1.11 3.44 1.175 3.405 1.175  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 3.89 0.31 4.01 0.31 4.01 0.605 3.89 0.605  ;
        POLYGON 3.89 0.8 4.01 0.8 4.01 1.235 3.89 1.235  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 2.375 0.26 2.41 0.26 2.41 0.085 1.445 0.085 1.445 0.45 1.38 0.45 1.38 0.085 0.675 0.085 0.675 0.36 0.61 0.36 0.61 0.085 0.3 0.085 0.3 0.28 0.235 0.28 0.235 0.085 0 0.085 0 -0.085 4.56 -0.085 4.56 0.085 4.195 0.085 4.195 0.34 4.13 0.34 4.13 0.085 3.59 0.085 3.59 0.395 3.525 0.395 3.525 0.085 2.475 0.085 2.475 0.26 2.51 0.26 2.51 0.325 2.375 0.325  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.615 0.62 0.715 0.62 0.715 0.755 0.615 0.755  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.18 0.61 0.315 0.61 0.315 0.745 0.18 0.745  ;
    END
  END CK
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.25 0.115 0.25 0.115 0.285 0.15 0.285 0.15 0.445 0.325 0.445 0.325 0.41 0.39 0.41 0.39 0.545 0.325 0.545 0.325 0.51 0.115 0.51 0.115 1.045 0.05 1.045  ;
        POLYGON 2.925 1.095 2.995 1.095 2.995 0.935 3.73 0.935 3.73 0.735 3.585 0.735 3.585 0.525 3.125 0.525 3.125 0.375 2.64 0.375 2.64 0.455 2.42 0.455 2.42 0.59 2.455 0.59 2.455 0.655 2.32 0.655 2.32 0.59 2.355 0.59 2.355 0.39 2.575 0.39 2.575 0.31 3.19 0.31 3.19 0.46 3.65 0.46 3.65 0.67 4.19 0.67 4.19 0.635 4.255 0.635 4.255 0.77 4.19 0.77 4.19 0.735 3.795 0.735 3.795 1.21 3.73 1.21 3.73 1 3.06 1 3.06 1.16 2.925 1.16  ;
        POLYGON 0.455 0.25 0.52 0.25 0.52 0.82 0.86 0.82 0.86 0.525 1.04 0.525 1.04 0.49 1.105 0.49 1.105 0.625 1.04 0.625 1.04 0.59 0.925 0.59 0.925 0.92 0.86 0.92 0.86 0.885 0.52 0.885 0.52 0.955 0.455 0.955  ;
        POLYGON 1.3 0.88 1.435 0.88 1.435 0.915 1.665 0.915 1.665 0.88 1.73 0.88 1.73 1.015 1.665 1.015 1.665 0.98 1.335 0.98 1.335 0.945 1.3 0.945  ;
        POLYGON 1.3 0.525 1.51 0.525 1.51 0.365 1.91 0.365 1.91 0.33 1.975 0.33 1.975 0.465 1.91 0.465 1.91 0.43 1.575 0.43 1.575 0.59 1.3 0.59  ;
        POLYGON 2.065 0.395 2.225 0.395 2.225 0.255 2.29 0.255 2.29 0.53 2.13 0.53 2.13 0.565 2.065 0.565  ;
        POLYGON 2.055 0.98 2.815 0.98 2.815 0.87 2.78 0.87 2.78 0.805 3.32 0.805 3.32 0.87 2.88 0.87 2.88 1.045 2.345 1.045 2.345 1.115 2.28 1.115 2.28 1.08 2.055 1.08  ;
        POLYGON 0.985 0.945 1.05 0.945 1.05 1.015 1.17 1.015 1.17 0.39 1.05 0.39 1.05 0.425 0.985 0.425 0.985 0.29 1.05 0.29 1.05 0.325 1.235 0.325 1.235 0.75 1.895 0.75 1.895 0.85 2.65 0.85 2.65 0.675 3.52 0.675 3.52 0.74 2.715 0.74 2.715 0.915 1.795 0.915 1.795 0.815 1.235 0.815 1.235 1.08 1.05 1.08 1.05 1.22 0.985 1.22  ;
  END
END DFFS_X2

MACRO DFFR_X1
  CLASS core ;
  FOREIGN DFFR_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 4.37 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 3.696 0.225 3.796 0.225 3.796 1.06 3.696 1.06  ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.511 0.405 2.181 0.405 2.181 0.375 2.411 0.375 2.411 0.2 2.515 0.2 2.515 0.16 2.615 0.16 2.615 0.2 3.056 0.2 3.056 0.485 3.301 0.485 3.301 0.55 2.991 0.55 2.991 0.265 2.476 0.265 2.476 0.44 2.236 0.44 2.236 0.47 1.511 0.47  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0.686 1.315 1.436 1.315 1.436 0.985 1.501 0.985 1.501 1.315 2.266 1.315 2.266 0.935 2.331 0.935 2.331 1.315 3.101 1.315 3.101 1.045 3.166 1.045 3.166 1.315 3.511 1.315 3.511 0.985 3.576 0.985 3.576 1.315 3.881 1.315 3.881 0.985 3.946 0.985 3.946 1.315 4.37 1.315 4.37 1.485 0 1.485 0 1.315 0.236 1.315 0.236 0.825 0.301 0.825 0.301 1.315 0.621 1.315 0.621 1.085 0.586 1.085 0.586 1.02 0.721 1.02 0.721 1.085 0.686 1.085  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 4.036 0.225 4.136 0.225 4.136 1.06 4.036 1.06  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 2.211 0.245 2.246 0.245 2.246 0.085 1.691 0.085 1.691 0.245 1.726 0.245 1.726 0.31 1.591 0.31 1.591 0.245 1.626 0.245 1.626 0.085 0.686 0.085 0.686 0.245 0.721 0.245 0.721 0.31 0.586 0.31 0.586 0.245 0.621 0.245 0.621 0.085 0.301 0.085 0.301 0.345 0.236 0.345 0.236 0.085 0 0.085 0 -0.085 4.37 -0.085 4.37 0.085 3.946 0.085 3.946 0.345 3.881 0.345 3.881 0.085 3.186 0.085 3.186 0.37 3.121 0.37 3.121 0.085 2.311 0.085 2.311 0.245 2.346 0.245 2.346 0.31 2.211 0.31  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.615 0.495 0.75 0.495 0.75 0.63 0.615 0.63  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.181 0.41 0.316 0.41 0.316 0.545 0.181 0.545  ;
    END
  END CK
  OBS
      LAYER M1 ;
        POLYGON 0.051 0.25 0.116 0.25 0.116 0.61 0.391 0.61 0.391 0.745 0.326 0.745 0.326 0.675 0.116 0.675 0.116 1.045 0.051 1.045  ;
        POLYGON 2.661 0.755 2.696 0.755 2.696 0.525 2.606 0.525 2.606 0.56 2.541 0.56 2.541 0.425 2.606 0.425 2.606 0.46 2.761 0.46 2.761 0.755 2.796 0.755 2.796 0.82 2.661 0.82  ;
        POLYGON 2.641 0.885 2.861 0.885 2.861 0.395 2.671 0.395 2.671 0.33 2.926 0.33 2.926 0.615 3.406 0.615 3.406 0.545 3.471 0.545 3.471 0.68 2.926 0.68 2.926 0.95 2.706 0.95 2.706 1.16 2.641 1.16  ;
        POLYGON 2.991 0.745 3.566 0.745 3.566 0.425 3.496 0.425 3.496 0.15 3.561 0.15 3.561 0.29 3.631 0.29 3.631 0.81 3.371 0.81 3.371 1.125 3.306 1.125 3.306 0.81 2.991 0.81  ;
        POLYGON 0.456 0.25 0.521 0.25 0.521 0.695 0.861 0.695 0.861 0.66 0.926 0.66 0.926 0.795 0.861 0.795 0.861 0.76 0.521 0.76 0.521 0.905 0.456 0.905  ;
        POLYGON 0.861 0.205 1.256 0.205 1.256 0.79 1.191 0.79 1.191 0.27 0.926 0.27 0.926 0.595 0.861 0.595  ;
        POLYGON 1.321 0.535 2.026 0.535 2.026 0.6 1.321 0.6  ;
        POLYGON 1.901 0.205 1.966 0.205 1.966 0.24 2.061 0.24 2.061 0.205 2.126 0.205 2.126 0.34 2.061 0.34 2.061 0.305 1.966 0.305 1.966 0.34 1.901 0.34  ;
        POLYGON 1.946 0.925 2.126 0.925 2.126 1.185 1.981 1.185 1.981 0.99 1.946 0.99  ;
        POLYGON 0.991 0.335 1.126 0.335 1.126 0.855 1.571 0.855 1.571 0.865 1.816 0.865 1.816 0.795 2.221 0.795 2.221 0.86 1.881 0.86 1.881 1.07 1.816 1.07 1.816 0.93 1.536 0.93 1.536 0.92 1.126 0.92 1.126 1.06 0.991 1.06  ;
        POLYGON 1.701 0.665 2.531 0.665 2.531 0.63 2.596 0.63 2.596 0.765 2.531 0.765 2.531 0.73 1.701 0.73  ;
  END
END DFFR_X1

MACRO DFFR_X2
  CLASS core ;
  FOREIGN DFFR_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 4.37 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 3.696 0.315 3.796 0.315 3.796 1.205 3.696 1.205  ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.511 0.405 2.181 0.405 2.181 0.375 2.411 0.375 2.411 0.2 2.515 0.2 2.515 0.16 2.615 0.16 2.615 0.2 3.056 0.2 3.056 0.515 3.301 0.515 3.301 0.58 2.991 0.58 2.991 0.265 2.476 0.265 2.476 0.44 2.236 0.44 2.236 0.47 1.511 0.47  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0.686 1.315 1.436 1.315 1.436 0.985 1.501 0.985 1.501 1.315 2.266 1.315 2.266 0.935 2.331 0.935 2.331 1.315 3.101 1.315 3.101 1.075 3.166 1.075 3.166 1.315 3.511 1.315 3.511 0.985 3.576 0.985 3.576 1.315 3.881 1.315 3.881 0.985 3.946 0.985 3.946 1.315 4.37 1.315 4.37 1.485 0 1.485 0 1.315 0.236 1.315 0.236 0.825 0.301 0.825 0.301 1.315 0.621 1.315 0.621 1.085 0.586 1.085 0.586 1.02 0.721 1.02 0.721 1.085 0.686 1.085  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 4.036 0.315 4.136 0.315 4.136 1.205 4.036 1.205  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 2.211 0.245 2.246 0.245 2.246 0.085 1.691 0.085 1.691 0.245 1.726 0.245 1.726 0.31 1.591 0.31 1.591 0.245 1.626 0.245 1.626 0.085 0.686 0.085 0.686 0.245 0.721 0.245 0.721 0.31 0.586 0.31 0.586 0.245 0.621 0.245 0.621 0.085 0.301 0.085 0.301 0.345 0.236 0.345 0.236 0.085 0 0.085 0 -0.085 4.37 -0.085 4.37 0.085 3.946 0.085 3.946 0.345 3.881 0.345 3.881 0.085 3.186 0.085 3.186 0.4 3.121 0.4 3.121 0.085 2.311 0.085 2.311 0.245 2.346 0.245 2.346 0.31 2.211 0.31  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.615 0.495 0.75 0.495 0.75 0.63 0.615 0.63  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.181 0.41 0.316 0.41 0.316 0.545 0.181 0.545  ;
    END
  END CK
  OBS
      LAYER M1 ;
        POLYGON 0.051 0.25 0.116 0.25 0.116 0.61 0.391 0.61 0.391 0.745 0.326 0.745 0.326 0.675 0.116 0.675 0.116 1.045 0.051 1.045  ;
        POLYGON 2.661 0.755 2.696 0.755 2.696 0.525 2.606 0.525 2.606 0.56 2.541 0.56 2.541 0.425 2.606 0.425 2.606 0.46 2.761 0.46 2.761 0.755 2.796 0.755 2.796 0.82 2.661 0.82  ;
        POLYGON 2.641 0.885 2.861 0.885 2.861 0.395 2.671 0.395 2.671 0.33 2.926 0.33 2.926 0.645 3.406 0.645 3.406 0.575 3.471 0.575 3.471 0.71 2.926 0.71 2.926 0.95 2.706 0.95 2.706 1.16 2.641 1.16  ;
        POLYGON 2.991 0.775 3.566 0.775 3.566 0.455 3.496 0.455 3.496 0.18 3.561 0.18 3.561 0.32 3.631 0.32 3.631 0.84 3.371 0.84 3.371 1.155 3.306 1.155 3.306 0.84 2.991 0.84  ;
        POLYGON 0.456 0.25 0.521 0.25 0.521 0.695 0.861 0.695 0.861 0.66 0.926 0.66 0.926 0.795 0.861 0.795 0.861 0.76 0.521 0.76 0.521 0.905 0.456 0.905  ;
        POLYGON 0.861 0.205 1.256 0.205 1.256 0.79 1.191 0.79 1.191 0.27 0.926 0.27 0.926 0.595 0.861 0.595  ;
        POLYGON 1.321 0.535 2.026 0.535 2.026 0.6 1.321 0.6  ;
        POLYGON 1.901 0.205 1.966 0.205 1.966 0.24 2.061 0.24 2.061 0.205 2.126 0.205 2.126 0.34 2.061 0.34 2.061 0.305 1.966 0.305 1.966 0.34 1.901 0.34  ;
        POLYGON 1.946 0.925 2.126 0.925 2.126 1.185 1.981 1.185 1.981 0.99 1.946 0.99  ;
        POLYGON 0.991 0.335 1.126 0.335 1.126 0.855 1.571 0.855 1.571 0.865 1.816 0.865 1.816 0.795 2.221 0.795 2.221 0.86 1.881 0.86 1.881 1.07 1.816 1.07 1.816 0.93 1.536 0.93 1.536 0.92 1.126 0.92 1.126 1.06 0.991 1.06  ;
        POLYGON 1.701 0.665 2.531 0.665 2.531 0.63 2.596 0.63 2.596 0.765 2.531 0.765 2.531 0.73 1.701 0.73  ;
  END
END DFFR_X2

MACRO SDFFSRX1  #SDFFRS_X1
  CLASS core ;
  #FOREIGN SDFFRS_X1 0.0 0.0 ;
  FOREIGN SDFFSRX1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 7.41 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 7.21 0.42 7.325 0.42 7.325 0.98 7.21 0.98  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
	CAPACITANCE 0.007796 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 3.11 0.508 4.095 0.508 4.095 0.598 5.105 0.598 5.105 0.663 4.03 0.663 4.03 0.573 3.11 0.573  ;
    END
  END SN
  PIN SE
    DIRECTION INPUT ;
	CAPACITANCE 0.001270 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.08 1.14 0.215 1.14 0.215 1.24 0.08 1.24  ;
    END
  END SE
  PIN RN
    DIRECTION INPUT ;
	CAPACITANCE 0.005751 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 3.81 0.638 3.945 0.638 3.945 0.728 4.96 0.728 4.96 0.793 3.88 0.793 3.88 0.703 3.81 0.703  ;
    END
  END RN
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 3.93 1.315 4.44 1.315 4.44 1.148 4.575 1.148 4.575 1.315 5.485 1.315 5.485 1.038 5.55 1.038 5.55 1.315 5.895 1.315 5.895 1.013 5.96 1.013 5.96 1.315 6.525 1.315 6.525 1.013 6.59 1.013 6.59 1.315 7.02 1.315 7.02 0.905 7.085 0.905 7.085 1.315 7.41 1.315 7.41 1.485 0 1.485 0 1.315 0.28 1.315 0.28 1.073 0.345 1.073 0.345 1.315 1.035 1.315 1.035 1.073 1.1 1.073 1.1 1.315 1.61 1.315 1.61 1.105 1.575 1.105 1.575 1.04 1.71 1.04 1.71 1.105 1.675 1.105 1.675 1.315 2.495 1.315 2.495 1.148 2.46 1.148 2.46 1.083 2.595 1.083 2.595 1.148 2.56 1.148 2.56 1.315 3.25 1.315 3.25 1.148 3.215 1.148 3.215 1.083 3.35 1.083 3.35 1.148 3.315 1.148 3.315 1.315 3.865 1.315 3.865 1.148 3.83 1.148 3.83 1.083 3.965 1.083 3.965 1.148 3.93 1.148  ;
    END
  END POWR  #VDD
  PIN Q
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 6.715 0.92 6.835 0.92 6.835 0.885 6.9 0.885 6.9 1.02 6.835 1.02 6.835 0.985 6.65 0.985 6.65 0.455 6.835 0.455 6.835 0.42 6.9 0.42 6.9 0.555 6.835 0.555 6.835 0.52 6.715 0.52  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
	CAPACITANCE 0.002952 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.325 0.368 0.425 0.368 0.425 0.3 0.525 0.3 0.525 0.368 0.975 0.368 0.975 0.513 1.01 0.513 1.01 0.578 0.875 0.578 0.875 0.433 0.325 0.433  ;
    END
  END SI
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 3.045 0.168 3.08 0.168 3.08 0.085 2.095 0.085 2.095 0.168 2.13 0.168 2.13 0.233 1.995 0.233 1.995 0.168 2.03 0.168 2.03 0.085 1.72 0.085 1.72 0.31 1.655 0.31 1.655 0.085 1.21 0.085 1.21 0.168 1.075 0.168 1.075 0.085 0.38 0.085 0.38 0.168 0.245 0.168 0.245 0.15 0.245 0.085 0 0.085 0 -0.085 7.41 -0.085 7.41 0.085 7.105 0.085 7.105 0.45 7.04 0.45 7.04 0.085 6.405 0.085 6.405 0.49 6.34 0.49 6.34 0.085 5.07 0.085 5.07 0.138 4.935 0.138 4.935 0.085 3.97 0.085 3.97 0.133 3.835 0.133 3.835 0.085 3.145 0.085 3.145 0.168 3.18 0.168 3.18 0.233 3.045 0.233  ;
    END
  END GRND  #VSS
  PIN D
    DIRECTION INPUT ;
	CAPACITANCE 0.002005 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.325 0.663 1 0.663 1 0.643 1.075 0.643 1.075 0.433 1.04 0.433 1.04 0.368 1.175 0.368 1.175 0.433 1.14 0.433 1.14 0.708 1.05 0.708 1.05 0.728 0.525 0.728 0.525 0.82 0.425 0.82 0.425 0.728 0.325 0.728  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
	CAPACITANCE 0.000397 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 1.555 0.44 1.69 0.44 1.69 0.54 1.555 0.54  ;
    END
  END CK
  OBS
      LAYER M1 ;
        POLYGON 0.04 0.823 0.075 0.823 0.075 0.173 0.14 0.173 0.14 0.498 0.81 0.498 0.81 0.563 0.14 0.563 0.14 0.823 0.175 0.823 0.175 0.888 0.04 0.888  ;
        POLYGON 3.245 0.178 3.54 0.178 3.54 0.243 3.245 0.243  ;
        POLYGON 2.92 0.638 3.405 0.638 3.405 0.733 3.61 0.733 3.61 0.698 3.745 0.698 3.745 0.763 3.71 0.763 3.71 0.798 3.305 0.798 3.305 0.703 2.92 0.703  ;
        POLYGON 1.87 1.063 2.33 1.063 2.33 0.903 2.725 0.903 2.725 1.063 3.085 1.063 3.085 0.863 3.735 0.863 3.735 0.858 4.435 0.858 4.435 0.923 3.76 0.923 3.76 0.928 3.15 0.928 3.15 1.128 2.66 1.128 2.66 0.968 2.395 0.968 2.395 1.128 1.87 1.128  ;
        POLYGON 4.475 0.338 4.51 0.338 4.51 0.243 4.235 0.243 4.235 0.178 4.575 0.178 4.575 0.338 4.61 0.338 4.61 0.403 4.475 0.403  ;
        POLYGON 5.135 0.893 5.17 0.893 5.17 0.533 4.16 0.533 4.16 0.413 2.69 0.413 2.69 0.578 1.84 0.578 1.84 0.38 1.805 0.38 1.805 0.315 2.015 0.315 2.015 0.513 2.625 0.513 2.625 0.413 2.59 0.413 2.59 0.348 4.225 0.348 4.225 0.468 5.235 0.468 5.235 0.893 5.27 0.893 5.27 0.958 5.135 0.958  ;
        POLYGON 4.97 1.053 5.005 1.053 5.005 0.958 4.565 0.958 4.565 1.083 4.03 1.083 4.03 1.018 4.5 1.018 4.5 0.893 5.07 0.893 5.07 1.053 5.335 1.053 5.335 0.438 5.4 0.438 5.4 1.118 4.97 1.118  ;
        POLYGON 4.675 0.338 4.71 0.338 4.71 0.303 5.735 0.303 5.735 0.828 6.025 0.828 6.025 0.793 6.09 0.793 6.09 1.153 6.395 1.153 6.395 0.685 6.46 0.685 6.46 1.218 6.025 1.218 6.025 0.893 5.735 0.893 5.735 0.978 5.67 0.978 5.67 0.368 4.81 0.368 4.81 0.403 4.675 0.403  ;
        POLYGON 5.965 0.41 6.03 0.41 6.03 0.555 6.52 0.555 6.52 0.52 6.585 0.52 6.585 0.655 6.52 0.655 6.52 0.62 6.22 0.62 6.22 1.088 6.155 1.088 6.155 0.62 5.965 0.62  ;
        POLYGON 6.78 0.685 6.845 0.685 6.845 0.72 7.08 0.72 7.08 0.685 7.145 0.685 7.145 0.82 6.78 0.82  ;
        POLYGON 1.23 0.903 1.525 0.903 1.525 0.968 1.23 0.968  ;
        POLYGON 1.78 0.903 2.075 0.903 2.075 0.968 1.78 0.968  ;
        POLYGON 0.625 0.823 1.1 0.823 1.1 0.773 1.24 0.773 1.24 0.303 0.965 0.303 0.965 0.273 0.625 0.273 0.625 0.208 1.02 0.208 1.02 0.238 1.305 0.238 1.305 0.773 2.235 0.773 2.235 0.808 2.27 0.808 2.27 0.873 2.135 0.873 2.135 0.838 1.165 0.838 1.165 0.888 0.625 0.888  ;
        POLYGON 2.46 0.153 2.525 0.153 2.525 0.448 2.46 0.448  ;
        POLYGON 1.49 0.643 2.855 0.643 2.855 0.998 2.79 0.998 2.79 0.708 1.37 0.708 1.37 0.315 1.525 0.315 1.525 0.38 1.49 0.38  ;
  END
END SDFFSRX1  #SDFFRS_X1

MACRO SDFFRS_X2
  CLASS core ;
  FOREIGN SDFFRS_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 7.41 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 7.21 0.42 7.325 0.42 7.325 0.98 7.21 0.98  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 3.11 0.508 4.105 0.508 4.105 0.6 5.115 0.6 5.115 0.665 4.04 0.665 4.04 0.573 3.11 0.573  ;
    END
  END SN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.08 1.14 0.215 1.14 0.215 1.24 0.08 1.24  ;
    END
  END SE
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 3.81 0.638 3.945 0.638 3.945 0.73 4.97 0.73 4.97 0.795 3.88 0.795 3.88 0.703 3.81 0.703  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 3.93 1.315 4.45 1.315 4.45 1.15 4.585 1.15 4.585 1.315 5.495 1.315 5.495 1.04 5.56 1.04 5.56 1.315 5.89 1.315 5.89 0.905 5.955 0.905 5.955 1.315 6.52 1.315 6.52 0.905 6.585 0.905 6.585 1.315 7.02 1.315 7.02 1.04 7.085 1.04 7.085 1.315 7.41 1.315 7.41 1.485 0 1.485 0 1.315 0.28 1.315 0.28 1.073 0.345 1.073 0.345 1.315 1.035 1.315 1.035 1.073 1.1 1.073 1.1 1.315 1.61 1.315 1.61 1.105 1.575 1.105 1.575 1.04 1.71 1.04 1.71 1.105 1.675 1.105 1.675 1.315 2.495 1.315 2.495 1.148 2.46 1.148 2.46 1.083 2.595 1.083 2.595 1.148 2.56 1.148 2.56 1.315 3.25 1.315 3.25 1.148 3.215 1.148 3.215 1.083 3.35 1.083 3.35 1.148 3.315 1.148 3.315 1.315 3.865 1.315 3.865 1.15 3.83 1.15 3.83 1.085 3.965 1.085 3.965 1.15 3.93 1.15  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 6.715 0.92 6.835 0.92 6.835 0.885 6.9 0.885 6.9 1.02 6.835 1.02 6.835 0.985 6.65 0.985 6.65 0.455 6.835 0.455 6.835 0.42 6.9 0.42 6.9 0.555 6.835 0.555 6.835 0.52 6.715 0.52  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.325 0.368 0.425 0.368 0.425 0.3 0.525 0.3 0.525 0.368 0.975 0.368 0.975 0.513 1.01 0.513 1.01 0.578 0.875 0.578 0.875 0.433 0.325 0.433  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 3.045 0.168 3.08 0.168 3.08 0.085 2.095 0.085 2.095 0.168 2.13 0.168 2.13 0.233 1.995 0.233 1.995 0.168 2.03 0.168 2.03 0.085 1.72 0.085 1.72 0.31 1.655 0.31 1.655 0.085 1.21 0.085 1.21 0.168 1.075 0.168 1.075 0.085 0.38 0.085 0.38 0.168 0.245 0.168 0.245 0.15 0.245 0.085 0 0.085 0 -0.085 7.41 -0.085 7.41 0.085 7.105 0.085 7.105 0.36 7.04 0.36 7.04 0.085 6.4 0.085 6.4 0.49 6.335 0.49 6.335 0.085 5.08 0.085 5.08 0.14 4.945 0.14 4.945 0.085 3.965 0.085 3.965 0.135 3.83 0.135 3.83 0.085 3.145 0.085 3.145 0.168 3.18 0.168 3.18 0.233 3.045 0.233  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.325 0.663 1 0.663 1 0.643 1.075 0.643 1.075 0.433 1.04 0.433 1.04 0.368 1.175 0.368 1.175 0.433 1.14 0.433 1.14 0.708 1.05 0.708 1.05 0.728 0.525 0.728 0.525 0.82 0.425 0.82 0.425 0.728 0.325 0.728  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.555 0.44 1.69 0.44 1.69 0.54 1.555 0.54  ;
    END
  END CK
  OBS
      LAYER M1 ;
        POLYGON 0.04 0.823 0.075 0.823 0.075 0.173 0.14 0.173 0.14 0.498 0.81 0.498 0.81 0.563 0.14 0.563 0.14 0.823 0.175 0.823 0.175 0.888 0.04 0.888  ;
        POLYGON 3.245 0.18 3.54 0.18 3.54 0.245 3.245 0.245  ;
        POLYGON 2.92 0.638 3.405 0.638 3.405 0.735 3.61 0.735 3.61 0.7 3.745 0.7 3.745 0.765 3.71 0.765 3.71 0.8 3.305 0.8 3.305 0.703 2.92 0.703  ;
        POLYGON 1.87 1.063 2.33 1.063 2.33 0.903 2.725 0.903 2.725 1.063 3.085 1.063 3.085 0.865 3.735 0.865 3.735 0.86 4.445 0.86 4.445 0.925 3.76 0.925 3.76 0.93 3.15 0.93 3.15 1.128 2.66 1.128 2.66 0.968 2.395 0.968 2.395 1.128 1.87 1.128  ;
        POLYGON 4.485 0.34 4.52 0.34 4.52 0.245 4.245 0.245 4.245 0.18 4.585 0.18 4.585 0.34 4.62 0.34 4.62 0.405 4.485 0.405  ;
        POLYGON 5.145 0.895 5.18 0.895 5.18 0.535 4.17 0.535 4.17 0.413 2.69 0.413 2.69 0.578 1.84 0.578 1.84 0.38 1.805 0.38 1.805 0.315 2.015 0.315 2.015 0.513 2.625 0.513 2.625 0.413 2.59 0.413 2.59 0.348 4.235 0.348 4.235 0.47 5.245 0.47 5.245 0.895 5.28 0.895 5.28 0.96 5.145 0.96  ;
        POLYGON 4.98 1.055 5.015 1.055 5.015 0.96 4.575 0.96 4.575 1.085 4.04 1.085 4.04 1.02 4.51 1.02 4.51 0.895 5.08 0.895 5.08 1.055 5.345 1.055 5.345 0.44 5.41 0.44 5.41 1.12 4.98 1.12  ;
        POLYGON 4.685 0.34 4.72 0.34 4.72 0.305 5.745 0.305 5.745 0.72 6.02 0.72 6.02 0.685 6.085 0.685 6.085 1.045 6.39 1.045 6.39 0.685 6.455 0.685 6.455 1.11 6.02 1.11 6.02 0.785 5.745 0.785 5.745 0.98 5.68 0.98 5.68 0.37 4.82 0.37 4.82 0.405 4.685 0.405  ;
        POLYGON 5.96 0.41 6.025 0.41 6.025 0.555 6.52 0.555 6.52 0.52 6.585 0.52 6.585 0.655 6.52 0.655 6.52 0.62 6.215 0.62 6.215 0.98 6.15 0.98 6.15 0.62 5.96 0.62  ;
        POLYGON 6.78 0.685 6.845 0.685 6.845 0.72 7.08 0.72 7.08 0.685 7.145 0.685 7.145 0.82 6.78 0.82  ;
        POLYGON 1.23 0.903 1.525 0.903 1.525 0.968 1.23 0.968  ;
        POLYGON 1.78 0.903 2.075 0.903 2.075 0.968 1.78 0.968  ;
        POLYGON 0.625 0.823 1.1 0.823 1.1 0.773 1.24 0.773 1.24 0.303 0.965 0.303 0.965 0.273 0.625 0.273 0.625 0.208 1.02 0.208 1.02 0.238 1.305 0.238 1.305 0.773 2.235 0.773 2.235 0.808 2.27 0.808 2.27 0.873 2.135 0.873 2.135 0.838 1.165 0.838 1.165 0.888 0.625 0.888  ;
        POLYGON 2.46 0.153 2.525 0.153 2.525 0.448 2.46 0.448  ;
        POLYGON 1.49 0.643 2.855 0.643 2.855 0.998 2.79 0.998 2.79 0.708 1.37 0.708 1.37 0.315 1.525 0.315 1.525 0.38 1.49 0.38  ;
  END
END SDFFRS_X2

MACRO TLATX1 #DLH_X1
  CLASS core ;
  FOREIGN TLATX1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 2.28 BY 1.4 ;
  PIN PWR
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.255 1.315 0.255 1.05 0.32 1.05 0.32 1.315 0.69 1.315 0.69 1.045 0.755 1.045 0.755 1.315 1.445 1.315 1.445 1.045 1.51 1.045 1.51 1.315 1.84 1.315 1.84 0.785 1.905 0.785 1.905 1.315 2.28 1.315 2.28 1.485 0 1.485  ;
    END
  END PWR
  PIN Q
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 2.01 0.415 2.11 0.415 2.11 0.775 2.01 0.775  ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 2.01 0.415 2.11 0.415 2.11 0.775 2.01 0.775  ;
    END
  END QN
  PIN GRND
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 2.28 -0.085 2.28 0.085 1.905 0.085 1.905 0.445 1.84 0.445 1.84 0.085 1.535 0.085 1.535 0.245 1.47 0.245 1.47 0.085 0.78 0.085 0.78 0.245 0.715 0.245 0.715 0.085 0.325 0.085 0.325 0.45 0.26 0.45 0.26 0.085 0 0.085  ;
    END
  END GRND
  PIN D
    DIRECTION INPUT ;
	CAPACITANCE 0.001178 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.555 0.15 0.62 0.15 0.62 0.31 0.835 0.31 0.835 0.44 0.905 0.44 0.905 0.54 0.835 0.54 0.835 0.85 0.77 0.85 0.77 0.375 0.555 0.375  ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
	CAPACITANCE 0.000734 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.2 0.745 0.335 0.745 0.335 0.88 0.2 0.88  ;
    END
  END C
  OBS
      LAYER M1 ;
        POLYGON 0.07 0.42 0.135 0.42 0.135 0.615 0.465 0.615 0.465 0.68 0.135 0.68 0.135 1.18 0.07 1.18  ;
        POLYGON 0.67 0.915 1.12 0.915 1.12 0.84 1.085 0.84 1.085 0.775 1.22 0.775 1.22 0.84 1.185 0.84 1.185 0.98 0.54 0.98 0.54 1.18 0.475 1.18 0.475 0.905 0.605 0.905 0.605 0.555 0.57 0.555 0.57 0.52 0.41 0.52 0.41 0.455 0.705 0.455 0.705 0.52 0.67 0.52  ;
        POLYGON 1.07 1.045 1.135 1.045 1.135 1.08 1.285 1.08 1.285 0.63 1.095 0.63 1.095 0.215 1.16 0.215 1.16 0.565 1.32 0.565 1.32 0.575 1.5 0.575 1.5 0.54 1.565 0.54 1.565 0.675 1.5 0.675 1.5 0.64 1.35 0.64 1.35 1.145 1.135 1.145 1.135 1.18 1.07 1.18  ;
        POLYGON 1.365 0.375 1.43 0.375 1.43 0.41 1.655 0.41 1.655 0.34 1.72 0.34 1.72 0.915 1.655 0.915 1.655 0.475 1.43 0.475 1.43 0.51 1.365 0.51  ;
  END
END TLATX1

MACRO DLH_X1
  CLASS core ;
  FOREIGN DLH_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 2.28 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.255 1.315 0.255 1.05 0.32 1.05 0.32 1.315 0.69 1.315 0.69 1.045 0.755 1.045 0.755 1.315 1.445 1.315 1.445 1.045 1.51 1.045 1.51 1.315 1.84 1.315 1.84 0.785 1.905 0.785 1.905 1.315 2.28 1.315 2.28 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 2.01 0.415 2.11 0.415 2.11 0.775 2.01 0.775  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 2.28 -0.085 2.28 0.085 1.905 0.085 1.905 0.445 1.84 0.445 1.84 0.085 1.535 0.085 1.535 0.245 1.47 0.245 1.47 0.085 0.78 0.085 0.78 0.245 0.715 0.245 0.715 0.085 0.325 0.085 0.325 0.45 0.26 0.45 0.26 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.555 0.15 0.62 0.15 0.62 0.31 0.835 0.31 0.835 0.44 0.905 0.44 0.905 0.54 0.835 0.54 0.835 0.85 0.77 0.85 0.77 0.375 0.555 0.375  ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.2 0.745 0.335 0.745 0.335 0.88 0.2 0.88  ;
    END
  END G
  OBS
      LAYER M1 ;
        POLYGON 0.07 0.42 0.135 0.42 0.135 0.615 0.465 0.615 0.465 0.68 0.135 0.68 0.135 1.18 0.07 1.18  ;
        POLYGON 0.67 0.915 1.12 0.915 1.12 0.84 1.085 0.84 1.085 0.775 1.22 0.775 1.22 0.84 1.185 0.84 1.185 0.98 0.54 0.98 0.54 1.18 0.475 1.18 0.475 0.905 0.605 0.905 0.605 0.555 0.57 0.555 0.57 0.52 0.41 0.52 0.41 0.455 0.705 0.455 0.705 0.52 0.67 0.52  ;
        POLYGON 1.07 1.045 1.135 1.045 1.135 1.08 1.285 1.08 1.285 0.63 1.095 0.63 1.095 0.215 1.16 0.215 1.16 0.565 1.32 0.565 1.32 0.575 1.5 0.575 1.5 0.54 1.565 0.54 1.565 0.675 1.5 0.675 1.5 0.64 1.35 0.64 1.35 1.145 1.135 1.145 1.135 1.18 1.07 1.18  ;
        POLYGON 1.365 0.375 1.43 0.375 1.43 0.41 1.655 0.41 1.655 0.34 1.72 0.34 1.72 0.915 1.655 0.915 1.655 0.475 1.43 0.475 1.43 0.51 1.365 0.51  ;
  END
END DLH_X1

MACRO DLH_X2
  CLASS core ;
  FOREIGN DLH_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 2.28 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.265 1.315 0.265 1.025 0.33 1.025 0.33 1.315 0.7 1.315 0.7 1.17 0.765 1.17 0.765 1.315 1.455 1.315 1.455 1.03 1.52 1.03 1.52 1.315 1.855 1.315 1.855 0.79 1.92 0.79 1.92 1.315 2.28 1.315 2.28 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 2.025 0.42 2.125 0.42 2.125 0.92 2.025 0.92  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 2.28 -0.085 2.28 0.085 1.935 0.085 1.935 0.45 1.87 0.45 1.87 0.085 1.585 0.085 1.585 0.255 1.52 0.255 1.52 0.085 0.83 0.085 0.83 0.255 0.765 0.255 0.765 0.085 0.33 0.085 0.33 0.425 0.265 0.425 0.265 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.605 0.15 0.67 0.15 0.67 0.32 0.845 0.32 0.845 0.44 0.905 0.44 0.905 0.54 0.845 0.54 0.845 0.86 0.78 0.86 0.78 0.385 0.605 0.385  ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.2 0.72 0.335 0.72 0.335 0.855 0.2 0.855  ;
    END
  END G
  OBS
      LAYER M1 ;
        POLYGON 0.035 0.395 0.145 0.395 0.145 0.59 0.45 0.59 0.45 0.655 0.135 0.655 0.135 1.155 0.035 1.155  ;
        POLYGON 0.68 0.925 1.13 0.925 1.13 0.825 1.095 0.825 1.095 0.76 1.23 0.76 1.23 0.825 1.195 0.825 1.195 0.99 0.54 0.99 0.54 1.2 0.475 1.2 0.475 0.925 0.615 0.925 0.615 0.53 0.495 0.53 0.495 0.495 0.42 0.495 0.42 0.43 0.555 0.43 0.555 0.465 0.715 0.465 0.715 0.53 0.68 0.53  ;
        POLYGON 1.08 1.055 1.145 1.055 1.145 1.09 1.295 1.09 1.295 0.62 1.145 0.62 1.145 0.225 1.21 0.225 1.21 0.555 1.36 0.555 1.36 0.62 1.51 0.62 1.51 0.585 1.575 0.585 1.575 0.72 1.51 0.72 1.51 0.685 1.36 0.685 1.36 1.155 1.145 1.155 1.145 1.19 1.08 1.19  ;
        POLYGON 1.415 0.385 1.48 0.385 1.48 0.42 1.685 0.42 1.685 0.385 1.785 0.385 1.785 0.92 1.67 0.92 1.67 0.52 1.415 0.52  ;
  END
END DLH_X2

MACRO DLL_X1
  CLASS core ;
  FOREIGN DLL_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 2.09 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.255 1.315 0.255 0.935 0.32 0.935 0.32 1.315 0.615 1.315 0.615 0.925 0.68 0.925 0.68 1.315 1.385 1.315 1.385 1.065 1.45 1.065 1.45 1.315 1.745 1.315 1.745 0.685 1.81 0.685 1.81 1.315 2.09 1.315 2.09 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.895 0.405 1.93 0.405 1.93 0.37 1.995 0.37 1.995 0.44 2.045 0.44 2.045 0.54 1.96 0.54 1.96 0.625 1.995 0.625 1.995 0.76 1.93 0.76 1.93 0.725 1.895 0.725  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0.235 0.32 0.27 0.32 0.27 0.085 0 0.085 0 -0.085 2.09 -0.085 2.09 0.085 1.79 0.085 1.79 0.49 1.725 0.49 1.725 0.085 1.45 0.085 1.45 0.505 1.385 0.505 1.385 0.085 0.68 0.085 0.68 0.415 0.615 0.415 0.615 0.085 0.335 0.085 0.335 0.32 0.37 0.32 0.37 0.455 0.235 0.455  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.615 0.545 0.715 0.545 0.715 0.68 0.615 0.68  ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.22 0.72 0.32 0.72 0.32 0.855 0.22 0.855  ;
    END
  END GN
  OBS
      LAYER M1 ;
        POLYGON 0.055 0.88 0.09 0.88 0.09 0.495 0.035 0.495 0.035 0.36 0.135 0.36 0.135 0.395 0.17 0.395 0.17 0.555 0.33 0.555 0.33 0.52 0.395 0.52 0.395 0.655 0.33 0.655 0.33 0.62 0.155 0.62 0.155 1.155 0.055 1.155  ;
        POLYGON 0.46 0.36 0.525 0.36 0.525 0.745 0.91 0.745 0.91 0.71 0.975 0.71 0.975 0.845 0.91 0.845 0.91 0.81 0.525 0.81 0.525 1.015 0.46 1.015  ;
        POLYGON 1.305 0.57 1.37 0.57 1.37 0.605 1.54 0.605 1.54 0.37 1.605 0.37 1.605 0.76 1.54 0.76 1.54 0.67 1.37 0.67 1.37 0.705 1.305 0.705  ;
        POLYGON 0.99 0.91 1.04 0.91 1.04 0.52 0.99 0.52 0.99 0.385 1.055 0.385 1.055 0.42 1.105 0.42 1.105 0.835 1.68 0.835 1.68 0.9 1.105 0.9 1.105 1.045 1.055 1.045 1.055 1.185 0.99 1.185  ;
  END
END DLL_X1

MACRO DLL_X2
  CLASS core ;
  FOREIGN DLL_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 2.09 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.255 1.315 0.255 0.935 0.32 0.935 0.32 1.315 0.615 1.315 0.615 0.93 0.68 0.93 0.68 1.315 1.385 1.315 1.385 0.965 1.45 0.965 1.45 1.315 1.745 1.315 1.745 0.68 1.81 0.68 1.81 1.315 2.09 1.315 2.09 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 1.895 0.435 1.93 0.435 1.93 0.4 1.995 0.4 1.995 0.44 2.045 0.44 2.045 0.54 1.96 0.54 1.96 0.625 1.995 0.625 1.995 0.9 1.93 0.9 1.93 0.76 1.895 0.76  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0.225 0.295 0.26 0.295 0.26 0.085 0 0.085 0 -0.085 2.09 -0.085 2.09 0.085 1.81 0.085 1.81 0.43 1.745 0.43 1.745 0.085 1.45 0.085 1.45 0.485 1.385 0.485 1.385 0.085 0.68 0.085 0.68 0.395 0.615 0.395 0.615 0.085 0.325 0.085 0.325 0.295 0.36 0.295 0.36 0.36 0.225 0.36  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.615 0.545 0.715 0.545 0.715 0.68 0.615 0.68  ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.22 0.72 0.32 0.72 0.32 0.855 0.22 0.855  ;
    END
  END GN
  OBS
      LAYER M1 ;
        POLYGON 0.055 0.88 0.09 0.88 0.09 0.495 0.035 0.495 0.035 0.36 0.135 0.36 0.135 0.395 0.17 0.395 0.17 0.555 0.33 0.555 0.33 0.52 0.395 0.52 0.395 0.655 0.33 0.655 0.33 0.62 0.155 0.62 0.155 1.155 0.055 1.155  ;
        POLYGON 0.46 0.36 0.525 0.36 0.525 0.745 0.91 0.745 0.91 0.71 0.975 0.71 0.975 0.845 0.91 0.845 0.91 0.81 0.525 0.81 0.525 1.015 0.46 1.015  ;
        POLYGON 1.305 0.55 1.37 0.55 1.37 0.585 1.54 0.585 1.54 0.4 1.605 0.4 1.605 0.76 1.54 0.76 1.54 0.65 1.37 0.65 1.37 0.685 1.305 0.685  ;
        POLYGON 0.99 0.91 1.04 0.91 1.04 0.5 0.99 0.5 0.99 0.365 1.055 0.365 1.055 0.4 1.105 0.4 1.105 0.835 1.68 0.835 1.68 0.9 1.105 0.9 1.105 1.045 1.055 1.045 1.055 1.185 0.99 1.185  ;
  END
END DLL_X2

MACRO DFFX1  #DFF_X1
  CLASS core ;
  #FOREIGN DFF_X1 0.0 0.0 ;
  FOREIGN DFFX1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 3.61 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 3.015 0.42 3.115 0.42 3.115 1.11 3.015 1.11  ;
    END
  END QN
  PIN POWR  #VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 2.63 1.315 3.31 1.315 3.31 1.035 3.375 1.035 3.375 1.315 3.61 1.315 3.61 1.485 0 1.485 0 1.315 0.235 1.315 0.235 0.84 0.3 0.84 0.3 1.315 0.94 1.315 0.94 1.025 1.005 1.025 1.005 1.315 1.81 1.315 1.81 0.99 1.875 0.99 1.875 1.315 2.565 1.315 2.565 1.125 2.53 1.125 2.53 1.025 2.665 1.025 2.665 1.125 2.63 1.125  ;
    END
  END POWR  #VDD
  PIN Q
    DIRECTION OUTPUT ;
	CAPACITANCE 0.008000 ;
    RESISTANCE 240.0 ;
    PORT
      LAYER M1 ;
        POLYGON 3.46 0.42 3.56 0.42 3.56 1.11 3.46 1.11  ;
    END
  END Q
  PIN GRND  #VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 2.53 0.225 2.565 0.225 2.565 0.085 1.87 0.085 1.87 0.225 1.905 0.225 1.905 0.29 1.77 0.29 1.77 0.225 1.805 0.225 1.805 0.085 1.005 0.085 1.005 0.325 0.94 0.325 0.94 0.085 0.3 0.085 0.3 0.245 0.235 0.245 0.235 0.085 0 0.085 0 -0.085 3.61 -0.085 3.61 0.085 3.3 0.085 3.3 0.54 3.235 0.54 3.235 0.085 2.63 0.085 2.63 0.225 2.665 0.225 2.665 0.29 2.53 0.29  ;
    END
  END GRND  #VSS
  PIN D
    DIRECTION INPUT ;
	CAPACITANCE 0.000705 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.985 0.65 1.085 0.65 1.085 0.785 0.985 0.785  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
	CAPACITANCE 0.000634 ;
    RESISTANCE 0.0 ;
    PORT
      LAYER M1 ;
        POLYGON 0.18 0.575 0.315 0.575 0.315 0.71 0.18 0.71  ;
    END
  END CK
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.215 0.115 0.215 0.115 0.41 0.29 0.41 0.29 0.375 0.355 0.375 0.355 0.51 0.29 0.51 0.29 0.475 0.115 0.475 0.115 1.01 0.05 1.01  ;
        POLYGON 2.19 0.85 2.795 0.85 2.795 1.175 3.18 1.175 3.18 0.815 3.245 0.815 3.245 1.24 2.73 1.24 2.73 0.915 2.255 0.915 2.255 1.11 2.19 1.11  ;
        POLYGON 0.42 0.165 0.875 0.165 0.875 0.39 1.535 0.39 1.535 0.525 1.47 0.525 1.47 0.455 0.81 0.455 0.81 0.23 0.555 0.23 0.555 0.87 0.42 0.87  ;
        POLYGON 0.645 0.295 0.745 0.295 0.745 0.52 1.405 0.52 1.405 0.59 1.8 0.59 1.8 0.655 1.34 0.655 1.34 0.585 0.745 0.585 0.745 1.145 0.645 1.145  ;
        POLYGON 1.43 0.19 1.495 0.19 1.495 0.225 1.705 0.225 1.705 0.425 1.99 0.425 1.99 0.49 1.64 0.49 1.64 0.29 1.495 0.29 1.495 0.325 1.43 0.325  ;
        POLYGON 0.815 0.85 1.485 0.85 1.485 1.01 1.68 1.01 1.68 0.85 1.99 0.85 1.99 0.915 1.745 0.915 1.745 1.075 1.485 1.075 1.485 1.11 1.42 1.11 1.42 0.915 0.88 0.915 0.88 0.985 0.815 0.985  ;
        POLYGON 1.18 0.65 1.245 0.65 1.245 0.685 1.28 0.685 1.28 0.72 2.065 0.72 2.065 0.425 2.27 0.425 2.27 0.39 2.335 0.39 2.335 0.525 2.27 0.525 2.27 0.49 2.13 0.49 2.13 0.82 2.065 0.82 2.065 0.785 1.615 0.785 1.615 0.945 1.55 0.945 1.55 0.785 1.18 0.785  ;
        POLYGON 2.19 0.19 2.255 0.19 2.255 0.225 2.465 0.225 2.465 0.55 2.795 0.55 2.795 0.615 2.4 0.615 2.4 0.29 2.255 0.29 2.255 0.325 2.19 0.325  ;
        POLYGON 2.45 0.68 2.86 0.68 2.86 0.295 2.925 0.295 2.925 1.11 2.86 1.11 2.86 0.745 2.45 0.745  ;
  END
END DFFX1  #DFF_X1

MACRO DFF_X2
  CLASS core ;
  FOREIGN DFF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 3.61 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 3.015 0.42 3.115 0.42 3.115 1.11 3.015 1.11  ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 2.63 1.315 3.31 1.315 3.31 1.17 3.375 1.17 3.375 1.315 3.61 1.315 3.61 1.485 0 1.485 0 1.315 0.235 1.315 0.235 0.84 0.3 0.84 0.3 1.315 0.94 1.315 0.94 1.025 1.005 1.025 1.005 1.315 1.81 1.315 1.81 0.99 1.875 0.99 1.875 1.315 2.565 1.315 2.565 1.125 2.53 1.125 2.53 1.025 2.665 1.025 2.665 1.125 2.63 1.125  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 3.46 0.42 3.56 0.42 3.56 1.11 3.46 1.11  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 2.53 0.225 2.565 0.225 2.565 0.085 1.87 0.085 1.87 0.225 1.905 0.225 1.905 0.29 1.77 0.29 1.77 0.225 1.805 0.225 1.805 0.085 1.005 0.085 1.005 0.325 0.94 0.325 0.94 0.085 0.3 0.085 0.3 0.245 0.235 0.245 0.235 0.085 0 0.085 0 -0.085 3.61 -0.085 3.61 0.085 3.37 0.085 3.37 0.45 3.305 0.45 3.305 0.085 2.63 0.085 2.63 0.225 2.665 0.225 2.665 0.29 2.53 0.29  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.985 0.65 1.085 0.65 1.085 0.785 0.985 0.785  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.18 0.575 0.315 0.575 0.315 0.71 0.18 0.71  ;
    END
  END CK
  OBS
      LAYER M1 ;
        POLYGON 0.05 0.215 0.115 0.215 0.115 0.41 0.29 0.41 0.29 0.375 0.355 0.375 0.355 0.51 0.29 0.51 0.29 0.475 0.115 0.475 0.115 1.01 0.05 1.01  ;
        POLYGON 2.19 0.85 2.795 0.85 2.795 1.175 3.18 1.175 3.18 0.815 3.245 0.815 3.245 1.24 2.73 1.24 2.73 0.915 2.255 0.915 2.255 1.11 2.19 1.11  ;
        POLYGON 0.42 0.165 0.875 0.165 0.875 0.39 1.535 0.39 1.535 0.525 1.47 0.525 1.47 0.455 0.81 0.455 0.81 0.23 0.555 0.23 0.555 0.87 0.42 0.87  ;
        POLYGON 0.645 0.295 0.745 0.295 0.745 0.52 1.405 0.52 1.405 0.59 1.8 0.59 1.8 0.655 1.34 0.655 1.34 0.585 0.745 0.585 0.745 1.145 0.645 1.145  ;
        POLYGON 1.43 0.19 1.495 0.19 1.495 0.225 1.705 0.225 1.705 0.425 1.99 0.425 1.99 0.49 1.64 0.49 1.64 0.29 1.495 0.29 1.495 0.325 1.43 0.325  ;
        POLYGON 0.815 0.85 1.485 0.85 1.485 1.01 1.68 1.01 1.68 0.85 1.99 0.85 1.99 0.915 1.745 0.915 1.745 1.075 1.485 1.075 1.485 1.11 1.42 1.11 1.42 0.915 0.88 0.915 0.88 0.985 0.815 0.985  ;
        POLYGON 1.18 0.65 1.245 0.65 1.245 0.685 1.28 0.685 1.28 0.72 2.065 0.72 2.065 0.425 2.27 0.425 2.27 0.39 2.335 0.39 2.335 0.525 2.27 0.525 2.27 0.49 2.13 0.49 2.13 0.82 2.065 0.82 2.065 0.785 1.615 0.785 1.615 0.945 1.55 0.945 1.55 0.785 1.18 0.785  ;
        POLYGON 2.19 0.19 2.255 0.19 2.255 0.225 2.465 0.225 2.465 0.55 2.795 0.55 2.795 0.615 2.4 0.615 2.4 0.29 2.255 0.29 2.255 0.325 2.19 0.325  ;
        POLYGON 2.45 0.68 2.86 0.68 2.86 0.295 2.925 0.295 2.925 1.11 2.86 1.11 2.86 0.745 2.45 0.745  ;
  END
END DFF_X2

MACRO SDFF_X1
  CLASS core ;
  FOREIGN SDFF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 4.94 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.425 0.42 0.56 0.42 0.56 0.83 0.425 0.83  ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 4.075 0.62 4.175 0.62 4.175 0.755 4.075 0.755  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.27 1.315 0.27 0.755 0.335 0.755 0.335 1.315 0.87 1.315 0.87 0.985 0.935 0.985 0.935 1.315 1.665 1.315 1.665 1.085 1.73 1.085 1.73 1.315 2.315 1.315 2.315 1.15 2.38 1.15 2.38 1.315 3.15 1.315 3.15 1.15 3.215 1.15 3.215 1.315 3.625 1.315 3.625 1 3.69 1 3.69 1.315 4.38 1.315 4.38 1 4.445 1 4.445 1.315 4.94 1.315 4.94 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.42 0.15 0.42 0.15 0.83 0.05 0.83  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 3.76 0.49 4.225 0.49 4.225 0.44 4.325 0.44 4.325 0.455 4.365 0.455 4.365 0.59 4.3 0.59 4.3 0.555 3.825 0.555 3.825 0.675 3.76 0.675  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 4.94 -0.085 4.94 0.085 4.45 0.085 4.45 0.15 4.45 0.325 4.385 0.325 4.385 0.085 3.575 0.085 3.575 0.325 3.51 0.325 3.51 0.085 3.165 0.085 3.165 0.27 3.1 0.27 3.1 0.085 2.375 0.085 2.375 0.26 2.31 0.26 2.31 0.085 1.735 0.085 1.735 0.415 1.67 0.415 1.67 0.085 0.935 0.085 0.935 0.415 0.87 0.415 0.87 0.085 0.335 0.085 0.335 0.54 0.27 0.54 0.27 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 3.6 0.52 3.665 0.52 3.665 0.74 3.95 0.74 3.95 0.82 4.3 0.82 4.3 0.785 4.365 0.785 4.365 0.92 4.325 0.92 4.325 0.96 4.225 0.96 4.225 0.885 3.885 0.885 3.885 0.805 3.6 0.805  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 3.275 0.755 3.375 0.755 3.375 0.89 3.275 0.89  ;
    END
  END CK
  OBS
      LAYER M1 ;
        POLYGON 2.82 0.955 3.405 0.955 3.405 1.09 3.34 1.09 3.34 1.02 2.72 1.02 2.72 0.885 2.755 0.885 2.755 0.72 1.795 0.72 1.795 0.755 1.73 0.755 1.73 0.72 1.36 0.72 1.36 0.755 1.295 0.755 1.295 0.62 1.36 0.62 1.36 0.655 1.73 0.655 1.73 0.62 1.795 0.62 1.795 0.655 2.755 0.655 2.755 0.465 2.72 0.465 2.72 0.4 2.87 0.4 2.87 0.435 2.905 0.435 2.905 0.47 3.34 0.47 3.34 0.4 3.405 0.4 3.405 0.535 2.82 0.535  ;
        POLYGON 3.535 0.87 3.82 0.87 3.82 0.985 4 0.985 4 0.95 4.065 0.95 4.065 1.085 4 1.085 4 1.05 3.755 1.05 3.755 0.935 3.47 0.935 3.47 0.665 3.11 0.665 3.11 0.735 3.045 0.735 3.045 0.6 3.47 0.6 3.47 0.39 3.64 0.39 3.64 0.325 4 0.325 4 0.29 4.065 0.29 4.065 0.425 4 0.425 4 0.39 3.705 0.39 3.705 0.455 3.535 0.455  ;
        POLYGON 4.57 0.295 4.69 0.295 4.69 1.22 4.57 1.22  ;
        POLYGON 0.65 0.18 0.75 0.18 0.75 1.105 0.65 1.105  ;
        POLYGON 0.88 0.82 1.065 0.82 1.065 1.02 1.25 1.02 1.25 0.985 1.315 0.985 1.315 1.12 1.25 1.12 1.25 1.085 1 1.085 1 0.885 0.88 0.885 0.88 0.92 0.815 0.92 0.815 0.48 0.88 0.48 0.88 0.515 1.175 0.515 1.175 0.33 1.25 0.33 1.25 0.295 1.315 0.295 1.315 0.43 1.24 0.43 1.24 0.58 0.88 0.58  ;
        POLYGON 1.17 0.785 1.235 0.785 1.235 0.82 1.975 0.82 1.975 1.115 1.855 1.115 1.855 0.885 1.235 0.885 1.235 0.92 1.17 0.92  ;
        POLYGON 2.05 0.15 2.17 0.15 2.17 0.46 2.05 0.46  ;
        POLYGON 2.075 0.82 2.45 0.82 2.45 0.785 2.515 0.785 2.515 0.92 2.45 0.92 2.45 0.885 2.175 0.885 2.175 1.235 2.075 1.235  ;
        POLYGON 1.42 0.455 1.485 0.455 1.485 0.49 1.855 0.49 1.855 0.295 1.975 0.295 1.975 0.525 2.59 0.525 2.59 0.455 2.655 0.455 2.655 0.59 1.855 0.59 1.855 0.555 1.485 0.555 1.485 0.59 1.42 0.59  ;
        POLYGON 2.235 0.325 2.3 0.325 2.3 0.36 2.465 0.36 2.465 0.185 2.72 0.185 2.72 0.15 2.785 0.15 2.785 0.285 2.72 0.285 2.72 0.25 2.53 0.25 2.53 0.425 2.3 0.425 2.3 0.46 2.235 0.46  ;
        POLYGON 2.24 0.95 2.305 0.95 2.305 0.985 2.51 0.985 2.51 1.135 2.775 1.135 2.775 1.1 2.84 1.1 2.84 1.235 2.775 1.235 2.775 1.2 2.445 1.2 2.445 1.05 2.305 1.05 2.305 1.085 2.24 1.085  ;
  END
END SDFF_X1

MACRO SDFF_X2
  CLASS core ;
  FOREIGN SDFF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE Free_OMC_Si2_PDK45nm ;
  SIZE 4.94 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.425 0.42 0.56 0.42 0.56 0.97 0.425 0.97  ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 4.075 0.62 4.175 0.62 4.175 0.755 4.075 0.755  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 1.315 0.27 1.315 0.27 0.89 0.335 0.89 0.335 1.315 0.87 1.315 0.87 0.985 0.935 0.985 0.935 1.315 1.665 1.315 1.665 1.085 1.73 1.085 1.73 1.315 2.315 1.315 2.315 1.15 2.38 1.15 2.38 1.315 3.15 1.315 3.15 1.15 3.215 1.15 3.215 1.315 3.625 1.315 3.625 1 3.69 1 3.69 1.315 4.38 1.315 4.38 1 4.445 1 4.445 1.315 4.94 1.315 4.94 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
        POLYGON 0.05 0.42 0.185 0.42 0.185 0.83 0.05 0.83  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 3.76 0.49 4.225 0.49 4.225 0.44 4.325 0.44 4.325 0.455 4.365 0.455 4.365 0.59 4.3 0.59 4.3 0.555 3.825 0.555 3.825 0.675 3.76 0.675  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        POLYGON 0 -0.085 4.94 -0.085 4.94 0.085 4.45 0.085 4.45 0.15 4.45 0.325 4.385 0.325 4.385 0.085 3.575 0.085 3.575 0.325 3.51 0.325 3.51 0.085 3.165 0.085 3.165 0.27 3.1 0.27 3.1 0.085 2.375 0.085 2.375 0.26 2.31 0.26 2.31 0.085 1.735 0.085 1.735 0.415 1.67 0.415 1.67 0.085 0.935 0.085 0.935 0.415 0.87 0.415 0.87 0.085 0.335 0.085 0.335 0.45 0.27 0.45 0.27 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 3.6 0.52 3.665 0.52 3.665 0.74 3.95 0.74 3.95 0.82 4.3 0.82 4.3 0.785 4.365 0.785 4.365 0.92 4.325 0.92 4.325 0.96 4.225 0.96 4.225 0.885 3.885 0.885 3.885 0.805 3.6 0.805  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
        POLYGON 3.275 0.755 3.375 0.755 3.375 0.89 3.275 0.89  ;
    END
  END CK
  OBS
      LAYER M1 ;
        POLYGON 2.82 0.955 3.405 0.955 3.405 1.09 3.34 1.09 3.34 1.02 2.72 1.02 2.72 0.885 2.755 0.885 2.755 0.72 1.795 0.72 1.795 0.755 1.73 0.755 1.73 0.72 1.36 0.72 1.36 0.755 1.295 0.755 1.295 0.62 1.36 0.62 1.36 0.655 1.73 0.655 1.73 0.62 1.795 0.62 1.795 0.655 2.755 0.655 2.755 0.465 2.72 0.465 2.72 0.4 2.87 0.4 2.87 0.435 2.905 0.435 2.905 0.47 3.34 0.47 3.34 0.4 3.405 0.4 3.405 0.535 2.82 0.535  ;
        POLYGON 3.535 0.87 3.82 0.87 3.82 0.985 4 0.985 4 0.95 4.065 0.95 4.065 1.085 4 1.085 4 1.05 3.755 1.05 3.755 0.935 3.47 0.935 3.47 0.665 3.11 0.665 3.11 0.735 3.045 0.735 3.045 0.6 3.47 0.6 3.47 0.39 3.64 0.39 3.64 0.325 4 0.325 4 0.29 4.065 0.29 4.065 0.425 4 0.425 4 0.39 3.705 0.39 3.705 0.455 3.535 0.455  ;
        POLYGON 4.57 0.295 4.69 0.295 4.69 1.22 4.57 1.22  ;
        POLYGON 0.65 0.18 0.75 0.18 0.75 1.105 0.65 1.105  ;
        POLYGON 0.88 0.82 1.065 0.82 1.065 1.02 1.25 1.02 1.25 0.985 1.315 0.985 1.315 1.12 1.25 1.12 1.25 1.085 1 1.085 1 0.885 0.88 0.885 0.88 0.92 0.815 0.92 0.815 0.48 0.88 0.48 0.88 0.515 1.175 0.515 1.175 0.33 1.25 0.33 1.25 0.295 1.315 0.295 1.315 0.43 1.24 0.43 1.24 0.58 0.88 0.58  ;
        POLYGON 1.17 0.785 1.235 0.785 1.235 0.82 1.975 0.82 1.975 1.115 1.855 1.115 1.855 0.885 1.235 0.885 1.235 0.92 1.17 0.92  ;
        POLYGON 2.05 0.15 2.17 0.15 2.17 0.46 2.05 0.46  ;
        POLYGON 2.075 0.82 2.45 0.82 2.45 0.785 2.515 0.785 2.515 0.92 2.45 0.92 2.45 0.885 2.175 0.885 2.175 1.235 2.075 1.235  ;
        POLYGON 1.42 0.455 1.485 0.455 1.485 0.49 1.855 0.49 1.855 0.295 1.975 0.295 1.975 0.525 2.59 0.525 2.59 0.455 2.655 0.455 2.655 0.59 1.855 0.59 1.855 0.555 1.485 0.555 1.485 0.59 1.42 0.59  ;
        POLYGON 2.235 0.325 2.3 0.325 2.3 0.36 2.465 0.36 2.465 0.185 2.72 0.185 2.72 0.15 2.785 0.15 2.785 0.285 2.72 0.285 2.72 0.25 2.53 0.25 2.53 0.425 2.3 0.425 2.3 0.46 2.235 0.46  ;
        POLYGON 2.24 0.95 2.305 0.95 2.305 0.985 2.51 0.985 2.51 1.135 2.775 1.135 2.775 1.1 2.84 1.1 2.84 1.235 2.775 1.235 2.775 1.2 2.445 1.2 2.445 1.05 2.305 1.05 2.305 1.085 2.24 1.085  ;
  END
END SDFF_X2

END LIBRARY
#
# End of file
#
