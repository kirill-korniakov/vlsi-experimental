VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.0025 ;

LAYER metal1
  TYPE ROUTING ;
  WIDTH 0.00034 ;
#  SPACING 0.065 ;
  PITCH 0.001 0.0007 ;
  DIRECTION HORIZONTAL ;
#  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.38 ;
#  THICKNESS 0.13 ;
  CAPACITANCE CPERSQDIST 20000.00 ;
  EDGECAPACITANCE 26.60 ;
END metal1

LAYER metal2
  TYPE ROUTING ;
  WIDTH 0.00037 ;
#  SPACING 0.07 ;
  PITCH 0.0001 0.0007 ;
  DIRECTION VERTICAL ;
#  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 259.00 ;
#  THICKNESS 0.14 ;
  CAPACITANCE CPERSQDIST 10000.00 ;
  EDGECAPACITANCE 23.15 ;
END metal2

LAYER metal3
  TYPE ROUTING ;
  WIDTH 0.00037 ;
#  SPACING 0.07 ;
  PITCH 0.001 0.0007 ;
  DIRECTION HORIZONTAL ;
#  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 259.00 ;
#  THICKNESS 0.14 ;
  CAPACITANCE CPERSQDIST 10000.00 ;
  EDGECAPACITANCE 23.15 ;
END metal3

SITE B5CSITE
#  SYMMETRY y ;
  CLASS core ;
  SIZE 0.001 BY 0.007 ;
END B5CSITE

MACRO AND2_X1
  ORIGIN 0 0 ;
  SITE B5CSITE ;
  SIZE 0.004 BY 0.007 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
  END VDD
  PIN A
    DIRECTION INPUT ;
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
  END VSS
  PIN B
    DIRECTION INPUT ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
  END Y
END AND2_X1

MACRO AND2_X2
  ORIGIN 0 0 ;
  SITE B5CSITE ;
  SIZE 0.004 BY 0.007 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
  END VDD
  PIN A
    DIRECTION INPUT ;
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
  END VSS
  PIN B
    DIRECTION INPUT ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
  END Y
END AND2_X2

MACRO AND2_X4
  ORIGIN 0 0 ;
  SITE B5CSITE ;
  SIZE 0.004 BY 0.007 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
  END VDD
  PIN A
    DIRECTION INPUT ;
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
  END VSS
  PIN B
    DIRECTION INPUT ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
  END Y
END AND2_X4

MACRO INV_X01
  ORIGIN 0 0 ;
  SITE B5CSITE ;
  SIZE 0.002 BY 0.007 ;
  PIN A
    DIRECTION INPUT ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
  END Y
END INV_X01

MACRO INV_X02
  ORIGIN 0 0 ;
  SITE B5CSITE ;
  SIZE 0.002 BY 0.007 ;
  PIN A
    DIRECTION INPUT ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
  END Y
END INV_X02

MACRO INV_X04
  ORIGIN 0 0 ;
  SITE B5CSITE ;
  SIZE 0.002 BY 0.007 ;
  PIN A
    DIRECTION INPUT ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
  END Y
END INV_X04

MACRO INV_X08
  ORIGIN 0 0 ;
  SITE B5CSITE ;
  SIZE 0.003 BY 0.007 ;
  PIN A
    DIRECTION INPUT ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
  END Y
END INV_X08

MACRO INV_X16
  ORIGIN 0 0 ;
  SITE B5CSITE ;
  SIZE 0.005 BY 0.007 ;
  PIN A
    DIRECTION INPUT ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
  END Y
END INV_X16

MACRO INV_X32
  ORIGIN 0 0 ;
  SITE B5CSITE ;
  SIZE 0.008 BY 0.007 ;
  PIN A
    DIRECTION INPUT ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
  END Y
END INV_X32

MACRO NAND2_X1
  ORIGIN 0 0 ;
  SITE B5CSITE ;
  SIZE 0.003 BY 0.007 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
  END VDD
  PIN A
    DIRECTION INPUT ;
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
  END VSS
  PIN B
    DIRECTION INPUT ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
  END Y
END NAND2_X1

MACRO NAND2_X2
  ORIGIN 0 0 ;
  SITE B5CSITE ;
  SIZE 0.003 BY 0.007 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
  END VDD
  PIN A
    DIRECTION INPUT ;
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
  END VSS
  PIN B
    DIRECTION INPUT ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
  END Y
END NAND2_X2

MACRO NAND2_X4
  ORIGIN 0 0 ;
  SITE B5CSITE ;
  SIZE 0.005 BY 0.007 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
  END VDD
  PIN A
    DIRECTION INPUT ;
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
  END VSS
  PIN B
    DIRECTION INPUT ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
  END Y
END NAND2_X4

MACRO OR2_X1
  ORIGIN 0 0 ;
  SITE B5CSITE ;
  SIZE 0.004 BY 0.007 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
  END VDD
  PIN A
    DIRECTION INPUT ;
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
  END VSS
  PIN B
    DIRECTION INPUT ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
  END Y
END OR2_X1

MACRO OR2_X2
  ORIGIN 0 0 ;
  SITE B5CSITE ;
  SIZE 0.004 BY 0.007 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
  END VDD
  PIN A
    DIRECTION INPUT ;
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
  END VSS
  PIN B
    DIRECTION INPUT ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
  END Y
END OR2_X2

MACRO OR2_X4
  ORIGIN 0 0 ;
  SITE B5CSITE ;
  SIZE 0.004 BY 0.007 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
  END VDD
  PIN A
    DIRECTION INPUT ;
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
  END VSS
  PIN B
    DIRECTION INPUT ;
  END B
  PIN Y
    DIRECTION OUTPUT ;
  END Y
END OR2_X4

END LIBRARY
#
# End of file
#
