#
#  180 nm Generic Library
#  Download from http://crete.cadence.com
#
# Export of the technology contained therein is governed by US Export
# Regulations. Diversion contrary to U.S. law is prohibited. Permission to make
# copies, either paper or electronic, of this work for personal or classroom use
# is granted without fee provided that the copies are not made or distributed for
# profit or commercial advantage. Users are free to use or modify content as
# appropriate as long as this notice appears in it. Information is provided 'as
# is' without warranty of any kind. No statement is made and no attempt has been
# made to examine the information, either with respect to operability, origin,
# authorship, or otherwise. Please use this information at your own risk. We
# recommend using it on a copy of your data to be sure you understand what it
# does under your conditions. Keep your master intact until you are satisfied
# with the use of this information within your environment. Please report any
# problems or enhancement requests to crete@cadence.com.  
# 
# Copyright 2003, Cadence Design Systems - All Rights Reserved
#
# LEF file generated by Abstract Generator version 5.5.13 on Apr  7 14:51:09 2005
#
# Contains LEF for all bins.
# Options:   [x] Antenna
#            [x] Geometry
#            [x] Technology

VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS

USEMINSPACING OBS ON ;
USEMINSPACING PIN OFF ;
CLEARANCEMEASURE EUCLIDEAN ;


MANUFACTURINGGRID 0.005 ;

LAYER Poly
  TYPE	MASTERSLICE ;
END Poly

LAYER Metal1
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		0.66  ;
  WIDTH		0.3 ;
  SPACING	0.3 ;
  SPACING	0.6 RANGE 10 100000  ;
  RESISTANCE	RPERSQ 0.101 ;
  CAPACITANCE	CPERSQDIST 0.00013153 ;
  EDGECAPACITANCE 8.770300e-05 ;
END Metal1

LAYER Via1
  TYPE	CUT ;
END Via1

LAYER Metal2
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		0.66  ;
  WIDTH		0.3 ;
  SPACING	0.3 ;
  SPACING	0.6 RANGE 10 100000  ;
  RESISTANCE	RPERSQ 0.101 ;
  CAPACITANCE	CPERSQDIST 7.0018e-05 ;
  EDGECAPACITANCE 8.311500e-05 ;
END Metal2

LAYER Via2
  TYPE	CUT ;
END Via2

LAYER Metal3
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		0.66  ;
  WIDTH		0.3 ;
  SPACING	0.3 ;
  SPACING	0.6 RANGE 10 100000  ;
  RESISTANCE	RPERSQ 0.101 ;
  CAPACITANCE	CPERSQDIST 6.3069e-05 ;
  EDGECAPACITANCE 1.002800e-04 ;
END Metal3

LAYER Via3
  TYPE	CUT ;
END Via3

LAYER Metal4
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		0.66  ;
  WIDTH		0.3 ;
  SPACING	0.3 ;
  SPACING	0.6 RANGE 10 100000  ;
  RESISTANCE	RPERSQ 0.101 ;
  CAPACITANCE	CPERSQDIST 5.3607e-05 ;
  EDGECAPACITANCE 8.298600e-05 ;
END Metal4

LAYER Via4
  TYPE	CUT ;
END Via4

LAYER Metal5
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		0.66  ;
  WIDTH		0.3 ;
  SPACING	0.3 ;
  SPACING	0.6 RANGE 10 100000  ;
  RESISTANCE	RPERSQ 0.045 ;
  CAPACITANCE	CPERSQDIST 3.144e-05 ;
  EDGECAPACITANCE 1.022400e-04 ;
END Metal5

LAYER Via5
  TYPE	CUT ;
END Via5

LAYER Metal6
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		0.66  ;
  WIDTH		0.3 ;
  SPACING	0.3 ;
  SPACING	0.6 RANGE 10 100000  ;
  RESISTANCE	RPERSQ 0.045 ;
  CAPACITANCE	CPERSQDIST 3.144e-05 ;
  EDGECAPACITANCE 1.022400e-04 ;
END Metal6

LAYER OVERLAP
  TYPE	OVERLAP ;
END OVERLAP

SPACING
  SAMENET Metal1  Metal1	0.300 ;
  SAMENET Metal2  Metal2	0.300  STACK ;
  SAMENET Metal3  Metal3	0.300  STACK ;
  SAMENET Metal4  Metal4	0.300  STACK ;
  SAMENET Metal5  Metal5	0.300  STACK ;
  SAMENET Metal6  Metal6	0.300 ;
  SAMENET Via1  Via1	0.300 ;
  SAMENET Via2  Via2	0.300 ;
  SAMENET Via3  Via3	0.300 ;
  SAMENET Via4  Via4	0.300 ;
  SAMENET Via1  Via2	0.000  STACK ;
  SAMENET Via2  Via3	0.000  STACK ;
  SAMENET Via3  Via4	0.000  STACK ;
  SAMENET Via4  Via5	0.000  STACK ;
END SPACING

VIA M2_M1 DEFAULT
  LAYER Metal1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER Via1 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER Metal2 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  RESISTANCE 6.400000e+00 ;
END M2_M1

VIA M3_M2 DEFAULT
  LAYER Metal2 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER Via2 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER Metal3 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  RESISTANCE 6.400000e+00 ;
END M3_M2

VIA M4_M3 DEFAULT
  LAYER Metal3 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER Via3 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER Metal4 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  RESISTANCE 6.400000e+00 ;
END M4_M3

VIA M5_M4 DEFAULT
  LAYER Metal4 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER Via4 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER Metal5 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  RESISTANCE 6.400000e+00 ;
END M5_M4

VIA M6_M5 DEFAULT
  LAYER Metal5 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER Via5 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER Metal6 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  RESISTANCE 6.400000e+00 ;
END M6_M5

VIA Via23_stack_north DEFAULT
  TOPOFSTACKONLY
  LAYER Metal2 ;
    RECT -0.200 -0.200 0.200 0.300 ;
  LAYER Via2 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER Metal3 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  RESISTANCE 6.400000e+00 ;
END Via23_stack_north

VIA Via23_stack_south DEFAULT
  TOPOFSTACKONLY
  LAYER Metal2 ;
    RECT -0.200 -0.300 0.200 0.200 ;
  LAYER Via2 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER Metal3 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  RESISTANCE 6.400000e+00 ;
END Via23_stack_south

VIA Via34_stack_east DEFAULT
  TOPOFSTACKONLY
  LAYER Metal3 ;
    RECT -0.200 -0.200 0.300 0.200 ;
  LAYER Via3 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER Metal4 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  RESISTANCE 6.400000e+00 ;
END Via34_stack_east

VIA Via34_stack_west DEFAULT
  TOPOFSTACKONLY
  LAYER Metal3 ;
    RECT -0.300 -0.200 0.200 0.200 ;
  LAYER Via3 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER Metal4 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  RESISTANCE 6.400000e+00 ;
END Via34_stack_west

VIA Via45_stack_north DEFAULT
  TOPOFSTACKONLY
  LAYER Metal4 ;
    RECT -0.200 -0.200 0.200 0.300 ;
  LAYER Via4 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER Metal5 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  RESISTANCE 2.540000e+00 ;
END Via45_stack_north

VIA Via45_stack_south DEFAULT
  TOPOFSTACKONLY
  LAYER Metal4 ;
    RECT -0.200 -0.300 0.200 0.200 ;
  LAYER Via4 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER Metal5 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  RESISTANCE 2.540000e+00 ;
END Via45_stack_south

VIA Via56_stack_east DEFAULT
  TOPOFSTACKONLY
  LAYER Metal5 ;
    RECT -0.200 -0.200 0.300 0.200 ;
  LAYER Via5 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER Metal6 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  RESISTANCE 2.540000e+00 ;
END Via56_stack_east

VIA Via56_stack_west DEFAULT
  TOPOFSTACKONLY
  LAYER Metal5 ;
    RECT -0.300 -0.200 0.200 0.200 ;
  LAYER Via5 ;
    RECT -0.100 -0.100 0.100 0.100 ;
  LAYER Metal6 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  RESISTANCE 2.540000e+00 ;
END Via56_stack_west


VIARULE Via12Array GENERATE
  LAYER Metal1 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.1 ;
    METALOVERHANG 0 ;
  LAYER Metal2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.1 ;
    METALOVERHANG 0 ;
  LAYER Via1 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.5 BY 0.5 ;
END Via12Array

VIARULE Via23Array GENERATE
  LAYER Metal3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.1 ;
    METALOVERHANG 0 ;
  LAYER Metal2 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.1 ;
    METALOVERHANG 0 ;
  LAYER Via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.5 BY 0.5 ;
END Via23Array

VIARULE Via34Array GENERATE
  LAYER Metal3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.1 ;
    METALOVERHANG 0 ;
  LAYER Metal4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.1 ;
    METALOVERHANG 0 ;
  LAYER Via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.5 BY 0.5 ;
END Via34Array

VIARULE Via45Array GENERATE
  LAYER Metal5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.1 ;
    METALOVERHANG 0 ;
  LAYER Metal4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.1 ;
    METALOVERHANG 0 ;
  LAYER Via4 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.5 BY 0.5 ;
END Via45Array

VIARULE Via56Array GENERATE
  LAYER Metal5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.1 ;
    METALOVERHANG 0 ;
  LAYER Metal6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.1 ;
    METALOVERHANG 0 ;
  LAYER Via5 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    SPACING 0.5 BY 0.5 ;
END Via56Array

VIARULE TURNMetal1 GENERATE
  LAYER Metal1 ;
    DIRECTION HORIZONTAL ;
  LAYER Metal1 ;
    DIRECTION VERTICAL ;
END TURNMetal1

VIARULE TURNMetal2 GENERATE
  LAYER Metal2 ;
    DIRECTION HORIZONTAL ;
  LAYER Metal2 ;
    DIRECTION VERTICAL ;
END TURNMetal2

VIARULE TURNMetal3 GENERATE
  LAYER Metal3 ;
    DIRECTION HORIZONTAL ;
  LAYER Metal3 ;
    DIRECTION VERTICAL ;
END TURNMetal3

VIARULE TURNMetal4 GENERATE
  LAYER Metal4 ;
    DIRECTION HORIZONTAL ;
  LAYER Metal4 ;
    DIRECTION VERTICAL ;
END TURNMetal4

VIARULE TURNMetal5 GENERATE
  LAYER Metal5 ;
    DIRECTION HORIZONTAL ;
  LAYER Metal5 ;
    DIRECTION VERTICAL ;
END TURNMetal5

VIARULE TURNMetal6 GENERATE
  LAYER Metal6 ;
    DIRECTION HORIZONTAL ;
  LAYER Metal6 ;
    DIRECTION VERTICAL ;
END TURNMetal6

SITE  CORE
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	0.660 BY 7.920 ;
END  CORE

MACRO TLATSRX1
  CLASS  CORE ;
  FOREIGN TLATSRX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.120 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.980 2.820 20.330 3.120 ;
        RECT 19.970 4.660 20.370 6.480 ;
        RECT 19.970 1.250 20.370 1.900 ;
        RECT 20.030 1.250 20.330 6.480 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 18.000 3.430 18.765 3.830 ;
        RECT 18.410 4.660 18.810 6.480 ;
        RECT 18.410 1.250 18.810 1.900 ;
        RECT 18.465 1.250 18.765 6.480 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.720 3.480 7.120 3.960 ;
        RECT 6.720 3.480 7.740 3.880 ;
    END
  END D
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.990 -0.540 5.890 0.650 ;
        RECT 0.000 -0.540 21.120 0.540 ;
        RECT 15.645 -0.540 19.590 0.650 ;
    END
  END GRND
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.600 3.480 6.000 3.960 ;
        RECT 5.600 3.480 6.420 3.780 ;
    END
  END G
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.400 2.820 12.290 3.120 ;
        RECT 13.350 2.690 13.750 3.090 ;
        RECT 11.790 2.690 13.750 2.990 ;
    END
  END RN
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 4.110 7.270 5.710 8.460 ;
        RECT 0.000 7.380 21.120 8.460 ;
        RECT 15.730 7.270 17.130 8.460 ;
    END
  END POWR
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.350 2.925 1.800 3.325 ;
        RECT 1.500 2.920 1.800 3.790 ;
    END
  END SN
  OBS 
      LAYER Metal1 ;
        RECT 0.650 1.390 1.150 1.790 ;
        RECT 0.650 4.660 1.150 5.460 ;
        RECT 0.650 1.390 0.950 6.820 ;
        RECT 0.650 6.420 1.050 6.820 ;
        RECT 1.530 4.660 1.930 6.880 ;
        RECT 1.530 1.150 1.930 1.790 ;
        RECT 4.110 4.660 4.510 6.770 ;
        RECT 4.110 1.150 4.510 1.790 ;
        RECT 3.225 3.560 3.625 4.060 ;
        RECT 3.225 3.760 5.110 4.060 ;
        RECT 4.810 3.760 5.110 5.460 ;
        RECT 4.810 4.660 5.290 5.460 ;
        RECT 6.490 4.660 6.890 6.880 ;
        RECT 6.490 1.040 6.890 1.790 ;
        RECT 7.270 1.140 7.850 1.790 ;
        RECT 2.555 1.390 3.110 1.790 ;
        RECT 4.320 2.695 8.030 2.995 ;
        RECT 7.630 2.695 8.030 3.115 ;
        RECT 2.555 2.960 4.620 3.260 ;
        RECT 2.555 1.390 2.855 5.260 ;
        RECT 2.510 4.660 2.910 5.260 ;
        RECT 4.890 1.390 5.290 1.790 ;
        RECT 4.890 1.390 5.190 2.395 ;
        RECT 9.030 1.790 9.430 2.190 ;
        RECT 3.385 2.095 9.330 2.395 ;
        RECT 3.225 2.195 3.625 2.595 ;
        RECT 9.830 5.080 10.230 6.880 ;
        RECT 11.255 1.040 11.655 1.540 ;
        RECT 12.690 4.960 13.090 6.880 ;
        RECT 12.690 1.040 13.090 1.790 ;
        RECT 9.030 3.295 9.430 3.795 ;
        RECT 14.250 3.130 14.650 3.795 ;
        RECT 9.030 3.495 14.650 3.795 ;
        RECT 10.365 2.090 14.650 2.390 ;
        RECT 14.250 2.090 14.650 2.590 ;
        RECT 10.365 2.090 10.765 2.820 ;
        RECT 16.030 4.660 16.430 6.770 ;
        RECT 8.230 1.140 10.475 1.440 ;
        RECT 14.430 1.140 14.830 1.790 ;
        RECT 9.730 1.140 10.475 1.540 ;
        RECT 8.230 1.140 8.630 1.790 ;
        RECT 14.430 1.490 15.730 1.790 ;
        RECT 9.730 1.140 10.030 2.995 ;
        RECT 8.330 2.695 10.030 2.995 ;
        RECT 16.030 3.860 16.430 4.260 ;
        RECT 15.430 3.960 16.430 4.260 ;
        RECT 8.330 4.360 15.730 4.660 ;
        RECT 11.140 4.360 11.440 6.480 ;
        RECT 15.430 1.490 15.730 5.265 ;
        RECT 14.430 4.965 15.730 5.265 ;
        RECT 8.330 2.695 8.630 6.480 ;
        RECT 8.230 4.660 8.630 6.480 ;
        RECT 11.090 5.080 11.490 6.480 ;
        RECT 14.430 4.960 14.830 6.780 ;
        RECT 16.030 1.150 16.430 2.190 ;
        RECT 16.810 1.790 17.210 2.190 ;
        RECT 16.910 2.590 17.610 2.990 ;
        RECT 16.910 1.790 17.210 5.460 ;
        RECT 16.810 4.660 17.210 5.460 ;
        RECT 19.190 4.660 19.590 6.880 ;
        RECT 19.190 1.150 19.590 1.900 ;
  END 
END TLATSRX1

MACRO TINVX1
  CLASS  CORE ;
  FOREIGN TINVX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.600 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN OE
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.320 3.240 1.720 3.830 ;
        RECT 1.320 3.430 1.850 3.830 ;
    END
  END OE
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.750 3.040 5.150 3.830 ;
        RECT 4.750 3.040 5.530 3.440 ;
    END
  END A
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.540 6.600 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.770 3.430 3.530 3.830 ;
        RECT 3.360 1.440 3.760 2.140 ;
        RECT 3.410 1.440 3.710 3.560 ;
        RECT 3.180 4.670 3.580 6.470 ;
        RECT 3.230 3.260 3.530 6.470 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 7.380 6.600 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.500 1.740 0.900 2.140 ;
        RECT 0.520 4.370 1.020 4.670 ;
        RECT 0.520 1.740 0.820 4.670 ;
        RECT 0.700 4.670 1.100 5.470 ;
        RECT 0.750 4.670 1.050 7.080 ;
        RECT 0.670 6.680 1.070 7.080 ;
        RECT 1.480 4.670 1.880 6.880 ;
        RECT 1.740 1.040 2.040 2.140 ;
        RECT 1.680 1.740 2.080 2.140 ;
        RECT 4.740 5.590 5.140 6.880 ;
        RECT 4.970 1.040 5.270 2.140 ;
        RECT 4.920 1.440 5.320 2.140 ;
        RECT 3.960 4.670 5.920 4.970 ;
        RECT 2.400 4.670 2.800 6.470 ;
        RECT 3.960 4.670 4.360 6.470 ;
        RECT 5.520 4.670 5.920 6.470 ;
        RECT 2.450 4.670 2.750 7.080 ;
        RECT 3.960 4.670 4.260 7.080 ;
        RECT 2.450 6.780 4.260 7.080 ;
        RECT 2.630 0.840 4.490 1.140 ;
        RECT 2.630 0.840 2.930 2.140 ;
        RECT 2.580 1.440 2.980 2.140 ;
        RECT 4.140 1.440 4.540 2.140 ;
        RECT 5.700 1.440 6.100 2.140 ;
        RECT 4.190 0.840 4.490 2.740 ;
        RECT 5.760 1.440 6.060 2.740 ;
        RECT 4.190 2.440 6.060 2.740 ;
  END 
END TINVX1

MACRO TLATX1
  CLASS  CORE ;
  FOREIGN TLATX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.220 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.890 1.290 10.190 6.320 ;
        RECT 9.890 3.480 10.380 3.780 ;
        RECT 9.820 4.520 10.220 6.320 ;
        RECT 9.820 1.290 10.220 1.940 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.260 1.290 7.660 1.940 ;
        RECT 7.360 4.520 7.760 6.340 ;
        RECT 7.360 2.820 7.740 3.120 ;
        RECT 7.360 1.290 7.660 4.220 ;
        RECT 7.280 3.920 7.580 4.980 ;
    END
  END QN
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.790 2.970 1.190 3.830 ;
        RECT 0.790 2.970 1.250 3.370 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.160 2.820 2.460 3.320 ;
        RECT 2.160 2.920 3.140 3.320 ;
    END
  END D
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.900 -0.540 7.800 0.650 ;
        RECT 0.000 -0.540 11.220 0.540 ;
    END
  END GRND
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.740 7.270 7.640 8.460 ;
        RECT 0.000 7.380 11.220 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 1.280 5.060 1.680 6.320 ;
        RECT 1.380 5.060 1.680 6.880 ;
        RECT 1.320 1.040 1.620 1.970 ;
        RECT 1.280 1.370 1.680 1.970 ;
        RECT 3.610 1.150 3.910 1.940 ;
        RECT 3.560 1.320 3.960 1.940 ;
        RECT 3.660 4.920 4.060 6.320 ;
        RECT 3.690 4.920 3.990 6.770 ;
        RECT 0.500 1.370 0.900 1.970 ;
        RECT 0.580 1.370 0.880 2.570 ;
        RECT 0.190 2.270 0.880 2.570 ;
        RECT 3.770 3.420 4.170 4.020 ;
        RECT 1.710 3.720 4.170 4.020 ;
        RECT 0.190 2.270 0.490 4.760 ;
        RECT 1.610 4.060 2.010 4.760 ;
        RECT 1.710 3.720 2.010 4.760 ;
        RECT 0.190 4.460 2.010 4.760 ;
        RECT 0.600 4.460 0.900 6.320 ;
        RECT 0.500 5.060 0.900 6.320 ;
        RECT 2.060 1.370 2.460 1.970 ;
        RECT 2.060 1.670 3.260 1.970 ;
        RECT 2.960 1.670 3.260 2.540 ;
        RECT 2.960 2.240 5.120 2.540 ;
        RECT 4.420 2.240 5.120 2.740 ;
        RECT 4.420 2.240 4.770 2.880 ;
        RECT 4.470 2.240 4.770 4.620 ;
        RECT 4.470 4.120 5.620 4.320 ;
        RECT 5.220 3.920 5.620 4.320 ;
        RECT 3.060 4.320 5.510 4.420 ;
        RECT 3.060 4.320 4.820 4.620 ;
        RECT 3.060 4.320 3.360 5.360 ;
        RECT 2.060 5.060 3.360 5.360 ;
        RECT 2.060 5.060 2.460 6.320 ;
        RECT 6.540 1.150 6.840 1.940 ;
        RECT 6.480 1.290 6.880 1.940 ;
        RECT 6.580 4.520 6.980 6.340 ;
        RECT 6.630 4.520 6.930 6.770 ;
        RECT 5.020 1.310 5.910 1.940 ;
        RECT 5.420 1.310 5.910 2.240 ;
        RECT 5.420 1.310 5.720 3.440 ;
        RECT 5.420 3.140 7.060 3.440 ;
        RECT 6.660 3.140 7.060 3.610 ;
        RECT 6.010 3.140 6.310 4.220 ;
        RECT 5.920 3.920 6.220 5.020 ;
        RECT 5.120 4.720 6.220 5.020 ;
        RECT 5.120 4.720 5.520 6.320 ;
        RECT 8.260 1.290 8.660 1.940 ;
        RECT 7.960 3.720 8.560 4.120 ;
        RECT 8.260 1.290 8.560 6.320 ;
        RECT 8.260 4.520 8.660 6.320 ;
        RECT 9.040 4.520 9.440 6.320 ;
        RECT 9.090 4.520 9.390 6.880 ;
        RECT 9.090 1.040 9.390 1.940 ;
        RECT 9.040 1.290 9.440 1.940 ;
  END 
END TLATX1

MACRO TBUFX4
  CLASS  CORE ;
  FOREIGN TBUFX4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.240 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN OE
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.760 2.820 3.160 3.290 ;
        RECT 2.760 2.890 3.280 3.290 ;
    END
  END OE
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.280 2.770 1.680 3.370 ;
        RECT 1.280 2.770 1.810 3.170 ;
    END
  END A
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 -0.540 3.430 0.650 ;
        RECT 8.060 -0.540 8.460 0.650 ;
        RECT 0.000 -0.540 9.240 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.940 4.250 5.240 6.670 ;
        RECT 8.180 1.440 8.580 2.370 ;
        RECT 6.500 2.680 8.480 2.980 ;
        RECT 8.180 1.440 8.480 2.980 ;
        RECT 6.620 1.440 7.020 2.370 ;
        RECT 6.620 1.440 6.920 2.980 ;
        RECT 6.400 4.850 6.800 6.670 ;
        RECT 6.500 2.670 6.800 6.670 ;
        RECT 4.940 4.250 6.800 4.550 ;
        RECT 6.070 3.430 6.800 3.830 ;
        RECT 4.840 4.850 5.240 6.670 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 4.160 7.270 8.080 8.460 ;
        RECT 0.000 7.380 9.240 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.500 4.360 0.900 6.880 ;
        RECT 1.280 1.880 2.680 2.180 ;
        RECT 1.280 1.250 1.680 2.250 ;
        RECT 2.280 1.250 2.680 2.250 ;
        RECT 3.060 4.360 3.460 6.880 ;
        RECT 3.130 1.150 3.430 2.250 ;
        RECT 3.060 1.250 3.460 2.250 ;
        RECT 4.060 4.850 4.460 6.670 ;
        RECT 4.160 4.850 4.460 6.770 ;
        RECT 4.060 1.040 4.460 3.040 ;
        RECT 0.500 1.250 0.900 2.250 ;
        RECT 0.500 1.250 0.800 4.060 ;
        RECT 0.500 3.760 4.630 4.060 ;
        RECT 2.290 3.760 2.590 7.080 ;
        RECT 4.230 3.760 4.630 4.450 ;
        RECT 1.280 4.420 2.680 4.720 ;
        RECT 1.280 4.360 1.680 7.080 ;
        RECT 2.280 4.360 2.680 7.080 ;
        RECT 5.620 4.850 6.020 6.670 ;
        RECT 5.670 4.850 5.970 6.770 ;
        RECT 7.180 4.850 7.580 6.670 ;
        RECT 7.230 4.850 7.530 6.770 ;
        RECT 5.890 0.840 7.760 1.140 ;
        RECT 5.890 0.840 6.190 2.370 ;
        RECT 7.460 0.840 7.760 2.370 ;
        RECT 4.840 1.640 6.240 1.940 ;
        RECT 5.840 1.440 6.240 2.370 ;
        RECT 7.400 1.440 7.800 2.370 ;
        RECT 4.840 0.840 5.240 3.040 ;
  END 
END TBUFX4

MACRO TBUFX8
  CLASS  CORE ;
  FOREIGN TBUFX8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.860 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN OE
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.520 3.380 5.200 3.780 ;
    END
  END OE
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 3.420 0.900 3.830 ;
        RECT 0.180 3.430 0.900 3.830 ;
    END
  END A
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 -0.540 3.300 0.650 ;
        RECT 12.500 -0.540 12.900 0.850 ;
        RECT 0.000 -0.540 13.860 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.060 3.960 7.360 6.670 ;
        RECT 11.640 4.560 12.040 6.670 ;
        RECT 11.690 3.960 11.990 6.670 ;
        RECT 7.060 3.960 11.990 4.260 ;
        RECT 11.080 1.450 11.480 2.950 ;
        RECT 9.570 3.250 11.430 3.550 ;
        RECT 11.130 1.450 11.430 3.550 ;
        RECT 10.700 3.250 11.100 4.260 ;
        RECT 10.080 4.560 10.480 6.670 ;
        RECT 10.130 3.960 10.430 6.670 ;
        RECT 9.520 1.450 9.920 2.950 ;
        RECT 9.570 1.450 9.870 3.550 ;
        RECT 8.520 4.560 8.920 6.670 ;
        RECT 8.570 3.960 8.870 6.670 ;
        RECT 6.960 4.560 7.360 6.670 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 7.270 11.680 8.460 ;
        RECT 0.000 7.380 13.860 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.500 4.880 0.900 6.670 ;
        RECT 0.600 4.880 0.900 6.770 ;
        RECT 2.060 4.880 2.460 6.670 ;
        RECT 2.100 4.880 2.400 6.770 ;
        RECT 2.890 1.150 3.190 2.610 ;
        RECT 2.840 1.550 3.240 2.610 ;
        RECT 3.620 4.880 4.020 6.670 ;
        RECT 3.680 4.880 3.980 6.770 ;
        RECT 0.550 0.950 2.410 1.250 ;
        RECT 0.550 0.950 0.850 2.610 ;
        RECT 0.500 1.550 0.900 2.610 ;
        RECT 2.060 1.550 2.460 2.610 ;
        RECT 3.620 1.550 4.020 2.610 ;
        RECT 2.110 0.950 2.410 3.240 ;
        RECT 3.670 1.550 3.970 3.240 ;
        RECT 2.110 2.940 3.970 3.240 ;
        RECT 5.180 4.880 5.580 6.670 ;
        RECT 5.210 4.880 5.510 6.770 ;
        RECT 5.400 1.040 5.800 2.340 ;
        RECT 6.180 4.560 6.580 6.670 ;
        RECT 6.230 4.560 6.530 6.770 ;
        RECT 1.280 1.550 1.680 2.610 ;
        RECT 6.180 3.760 6.580 4.160 ;
        RECT 5.580 3.860 6.580 4.160 ;
        RECT 5.580 3.860 5.880 4.580 ;
        RECT 1.330 4.280 5.880 4.580 ;
        RECT 1.330 1.550 1.630 6.670 ;
        RECT 2.890 4.280 3.190 6.670 ;
        RECT 4.470 4.280 4.770 6.670 ;
        RECT 1.280 4.880 1.680 6.670 ;
        RECT 2.840 4.880 3.240 6.670 ;
        RECT 4.400 4.880 4.800 6.670 ;
        RECT 6.960 1.040 7.360 2.340 ;
        RECT 7.740 4.560 8.140 6.670 ;
        RECT 7.790 4.560 8.090 6.770 ;
        RECT 9.300 4.560 9.700 6.670 ;
        RECT 9.370 4.560 9.670 6.770 ;
        RECT 10.860 4.560 11.260 6.670 ;
        RECT 10.910 4.560 11.210 6.770 ;
        RECT 7.740 0.850 12.200 1.150 ;
        RECT 8.790 0.850 9.090 2.950 ;
        RECT 10.360 0.850 10.660 2.950 ;
        RECT 11.900 0.850 12.200 2.950 ;
        RECT 4.620 0.840 5.020 2.340 ;
        RECT 6.180 0.840 6.580 2.340 ;
        RECT 7.740 0.840 8.140 2.340 ;
        RECT 4.690 0.840 4.990 2.940 ;
        RECT 6.230 0.840 6.530 2.940 ;
        RECT 7.790 0.840 8.090 2.940 ;
        RECT 4.690 2.640 8.090 2.940 ;
        RECT 8.740 1.450 9.140 2.950 ;
        RECT 10.300 1.450 10.700 2.950 ;
        RECT 11.860 1.450 12.260 2.950 ;
  END 
END TBUFX8

MACRO TBUFX1
  CLASS  CORE ;
  FOREIGN TBUFX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.940 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN OE
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.790 4.090 1.190 5.010 ;
        RECT 0.680 4.610 1.190 5.010 ;
    END
  END OE
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.080 3.940 2.510 4.340 ;
        RECT 2.110 3.940 2.510 4.490 ;
    END
  END A
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 -0.540 5.300 0.650 ;
        RECT 0.000 -0.540 5.940 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.840 1.250 5.240 1.900 ;
        RECT 4.840 4.850 5.240 6.670 ;
        RECT 4.940 1.250 5.240 6.670 ;
        RECT 4.800 2.820 5.240 3.120 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.530 7.270 5.170 8.460 ;
        RECT 0.000 7.380 5.940 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.500 5.410 0.900 6.670 ;
        RECT 0.530 5.410 0.830 6.770 ;
        RECT 0.550 1.150 0.850 1.650 ;
        RECT 0.500 1.250 0.900 1.650 ;
        RECT 1.280 1.250 1.680 2.640 ;
        RECT 1.280 2.240 2.210 2.640 ;
        RECT 1.810 2.240 2.210 3.380 ;
        RECT 2.310 1.150 2.610 1.900 ;
        RECT 2.280 1.250 2.680 1.900 ;
        RECT 3.060 5.410 3.460 6.670 ;
        RECT 3.110 5.410 3.410 6.770 ;
        RECT 4.060 4.850 4.460 6.670 ;
        RECT 4.100 4.850 4.400 6.770 ;
        RECT 3.060 1.320 4.460 1.620 ;
        RECT 3.060 1.250 3.460 1.900 ;
        RECT 4.060 1.250 4.460 1.900 ;
        RECT 2.590 2.980 2.990 3.380 ;
        RECT 2.590 3.080 4.230 3.380 ;
        RECT 3.930 3.080 4.230 4.550 ;
        RECT 3.930 4.040 4.630 4.440 ;
        RECT 3.460 4.250 4.620 4.550 ;
        RECT 3.460 4.250 3.760 5.110 ;
        RECT 2.380 4.810 3.760 5.110 ;
        RECT 1.280 5.480 2.680 5.780 ;
        RECT 1.280 5.410 1.680 6.670 ;
        RECT 2.380 4.810 2.680 6.670 ;
        RECT 2.280 5.410 2.680 6.670 ;
  END 
END TBUFX1

MACRO TBUFX2
  CLASS  CORE ;
  FOREIGN TBUFX2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.940 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN OE
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.970 2.560 1.370 3.140 ;
        RECT 0.970 2.740 3.590 3.140 ;
    END
  END OE
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.880 4.140 2.280 4.540 ;
        RECT 1.880 4.140 2.460 4.440 ;
    END
  END A
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 -0.540 2.100 0.650 ;
        RECT 0.000 -0.540 5.940 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.930 4.240 4.230 6.670 ;
        RECT 4.720 2.830 5.100 3.130 ;
        RECT 3.930 4.240 5.020 4.540 ;
        RECT 4.720 0.840 5.020 4.540 ;
        RECT 4.620 0.840 5.020 2.340 ;
        RECT 3.840 4.850 4.240 6.670 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.530 7.270 5.170 8.460 ;
        RECT 0.000 7.380 5.940 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.500 5.410 0.900 6.670 ;
        RECT 0.530 5.410 0.830 6.770 ;
        RECT 0.550 1.150 0.850 1.650 ;
        RECT 0.500 1.250 0.900 1.650 ;
        RECT 1.330 1.050 1.630 1.650 ;
        RECT 1.280 1.250 1.680 1.650 ;
        RECT 2.060 5.410 2.460 6.670 ;
        RECT 2.120 5.410 2.420 6.770 ;
        RECT 3.060 4.850 3.460 6.670 ;
        RECT 3.110 4.850 3.410 6.770 ;
        RECT 3.060 1.040 3.460 2.340 ;
        RECT 3.840 0.840 4.240 2.340 ;
        RECT 2.060 1.250 2.460 1.650 ;
        RECT 2.130 1.250 2.430 2.250 ;
        RECT 0.370 1.950 2.430 2.250 ;
        RECT 0.370 3.540 4.420 3.840 ;
        RECT 4.020 3.540 4.420 3.940 ;
        RECT 0.370 1.950 0.670 5.110 ;
        RECT 0.370 4.810 1.580 5.110 ;
        RECT 1.280 4.810 1.580 6.670 ;
        RECT 1.280 5.410 1.680 6.670 ;
        RECT 4.620 4.850 5.020 6.670 ;
        RECT 4.670 4.850 4.970 6.770 ;
  END 
END TBUFX2

MACRO FILL8
  CLASS  CORE ;
  FOREIGN FILL8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.540 -0.540 3.940 0.650 ;
        RECT 0.000 -0.540 5.280 0.540 ;
    END
  END GRND
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.930 7.260 3.330 8.460 ;
        RECT 0.000 7.380 5.280 8.460 ;
    END
  END POWR
END FILL8

MACRO ADDFX1
  CLASS  CORE ;
  FOREIGN ADDFX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.420 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.690 2.820 3.990 4.590 ;
        RECT 9.110 2.820 9.510 3.460 ;
        RECT 3.690 2.820 9.510 3.120 ;
        RECT 6.540 3.560 6.940 3.960 ;
        RECT 6.070 3.560 6.940 3.860 ;
        RECT 6.070 2.820 6.470 3.860 ;
        RECT 3.600 4.190 4.000 4.590 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.750 4.680 5.150 5.080 ;
        RECT 9.110 4.070 9.510 4.470 ;
        RECT 5.460 4.270 9.500 4.570 ;
        RECT 4.750 4.780 5.860 5.080 ;
        RECT 5.460 4.140 5.860 5.080 ;
    END
  END B
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 22.290 2.840 22.590 6.480 ;
        RECT 23.470 1.250 23.870 1.900 ;
        RECT 22.290 2.840 23.820 3.140 ;
        RECT 23.520 1.250 23.820 3.140 ;
        RECT 22.190 4.660 22.590 6.480 ;
    END
  END S
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.740 -0.540 1.440 0.650 ;
        RECT 10.600 -0.540 12.000 0.650 ;
        RECT 0.000 -0.540 24.420 0.540 ;
    END
  END GRND
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.440 3.430 8.510 3.830 ;
        RECT 8.110 3.430 8.510 3.970 ;
    END
  END CI
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.820 7.270 2.250 8.460 ;
        RECT 0.000 7.380 24.420 8.460 ;
        RECT 22.110 7.270 23.510 8.460 ;
        RECT 14.430 7.270 15.830 8.460 ;
    END
  END POWR
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 3.480 1.400 3.780 ;
        RECT 1.120 4.540 1.520 6.360 ;
        RECT 1.120 1.250 1.520 1.900 ;
        RECT 1.100 1.320 1.400 5.280 ;
    END
  END CO
  OBS 
      LAYER Metal1 ;
        RECT 1.900 4.540 2.300 6.360 ;
        RECT 1.950 4.540 2.250 6.770 ;
        RECT 1.940 1.040 2.240 1.900 ;
        RECT 1.900 1.250 2.300 1.900 ;
        RECT 3.680 5.490 4.080 6.750 ;
        RECT 3.680 0.920 4.480 1.320 ;
        RECT 4.460 5.490 4.860 6.750 ;
        RECT 4.510 5.490 4.810 6.880 ;
        RECT 4.860 1.040 5.260 1.320 ;
        RECT 5.460 5.490 5.860 6.750 ;
        RECT 5.510 5.490 5.810 6.880 ;
        RECT 5.860 1.040 6.260 1.320 ;
        RECT 7.240 5.490 7.640 6.750 ;
        RECT 7.330 5.490 7.630 6.880 ;
        RECT 7.640 1.040 8.040 1.320 ;
        RECT 6.290 4.890 8.370 5.190 ;
        RECT 6.290 4.890 6.590 6.750 ;
        RECT 8.070 4.890 8.370 6.750 ;
        RECT 6.240 5.490 6.640 6.750 ;
        RECT 8.020 5.490 8.420 6.750 ;
        RECT 6.640 0.920 7.040 1.320 ;
        RECT 8.420 0.920 9.220 1.320 ;
        RECT 6.740 0.920 7.040 1.920 ;
        RECT 8.500 0.920 8.800 1.920 ;
        RECT 6.740 1.620 8.800 1.920 ;
        RECT 10.560 5.210 10.960 6.470 ;
        RECT 10.590 5.210 10.890 6.880 ;
        RECT 11.020 1.150 11.320 2.140 ;
        RECT 11.010 1.740 11.410 2.140 ;
        RECT 2.900 0.920 3.300 1.320 ;
        RECT 9.600 0.920 10.250 1.320 ;
        RECT 2.900 2.220 10.250 2.520 ;
        RECT 9.950 2.860 12.530 3.160 ;
        RECT 12.130 2.800 12.530 3.200 ;
        RECT 1.820 3.730 2.220 4.130 ;
        RECT 1.820 3.830 3.200 4.130 ;
        RECT 2.900 0.920 3.200 6.750 ;
        RECT 9.950 0.920 10.250 5.950 ;
        RECT 8.800 5.650 10.250 5.950 ;
        RECT 2.900 5.490 3.300 6.750 ;
        RECT 8.800 5.490 9.200 6.750 ;
        RECT 13.040 3.460 13.440 3.860 ;
        RECT 10.620 3.560 13.440 3.860 ;
        RECT 10.620 3.480 11.020 3.880 ;
        RECT 15.300 5.210 15.700 6.470 ;
        RECT 15.350 5.210 15.650 6.770 ;
        RECT 15.410 1.040 15.710 1.850 ;
        RECT 15.350 1.450 15.750 1.850 ;
        RECT 14.630 4.610 16.600 4.910 ;
        RECT 14.550 4.620 14.850 6.470 ;
        RECT 11.340 5.210 11.740 6.470 ;
        RECT 13.820 5.920 14.920 6.220 ;
        RECT 12.340 4.870 12.740 6.470 ;
        RECT 11.340 6.170 12.740 6.470 ;
        RECT 14.520 5.210 14.920 6.470 ;
        RECT 16.400 4.620 16.700 6.470 ;
        RECT 16.300 5.210 16.700 6.470 ;
        RECT 12.410 4.870 12.710 7.070 ;
        RECT 13.830 5.920 14.130 7.070 ;
        RECT 12.410 6.770 14.130 7.070 ;
        RECT 12.850 0.840 14.910 1.140 ;
        RECT 16.770 0.840 17.170 1.240 ;
        RECT 12.850 0.840 13.150 1.950 ;
        RECT 14.570 1.450 14.970 1.850 ;
        RECT 12.790 1.450 13.190 1.950 ;
        RECT 11.790 1.650 13.190 1.950 ;
        RECT 11.790 1.650 12.190 2.140 ;
        RECT 14.610 0.840 14.910 2.460 ;
        RECT 16.820 0.840 17.120 2.460 ;
        RECT 14.610 2.160 17.120 2.460 ;
        RECT 17.080 5.210 17.480 6.470 ;
        RECT 17.130 5.210 17.430 6.880 ;
        RECT 17.550 1.040 17.950 1.240 ;
        RECT 18.080 4.870 18.480 6.470 ;
        RECT 18.140 4.870 18.440 6.880 ;
        RECT 18.550 1.040 18.950 1.340 ;
        RECT 18.860 4.870 19.260 6.470 ;
        RECT 17.420 2.240 17.820 2.690 ;
        RECT 19.460 2.270 19.860 2.690 ;
        RECT 17.420 2.390 19.860 2.690 ;
        RECT 19.640 4.870 20.040 6.470 ;
        RECT 19.330 0.840 20.130 1.340 ;
        RECT 14.430 3.290 14.830 3.690 ;
        RECT 19.990 3.300 20.390 3.700 ;
        RECT 14.440 3.400 20.390 3.700 ;
        RECT 20.510 0.840 21.310 1.340 ;
        RECT 21.410 4.660 21.810 6.480 ;
        RECT 21.470 4.660 21.770 6.770 ;
        RECT 21.470 4.660 21.610 6.880 ;
        RECT 21.690 0.840 22.090 1.340 ;
        RECT 13.570 1.450 14.070 1.950 ;
        RECT 21.690 0.840 21.990 1.950 ;
        RECT 20.710 1.650 21.990 1.950 ;
        RECT 13.770 4.000 21.990 4.300 ;
        RECT 21.590 3.860 21.990 4.300 ;
        RECT 13.770 1.450 14.070 4.560 ;
        RECT 13.180 4.260 14.070 4.560 ;
        RECT 13.180 4.260 13.480 6.470 ;
        RECT 13.120 4.870 13.520 6.470 ;
        RECT 20.710 1.650 21.010 6.470 ;
        RECT 20.420 4.870 21.010 6.470 ;
        RECT 22.820 1.040 23.120 1.680 ;
        RECT 22.690 1.250 23.090 1.900 ;
  END 
END ADDFX1

MACRO ADDHX1
  CLASS  CORE ;
  FOREIGN ADDHX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.160 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 10.690 4.080 11.090 4.810 ;
        RECT 10.520 4.410 11.090 4.810 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.470 2.650 7.870 3.050 ;
        RECT 9.270 1.390 9.780 1.790 ;
        RECT 7.470 2.750 9.570 3.050 ;
        RECT 9.270 1.360 9.570 3.050 ;
        RECT 8.050 2.750 8.450 3.210 ;
    END
  END B
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.060 0.840 2.460 2.240 ;
        RECT 3.880 2.770 4.490 3.170 ;
        RECT 2.330 3.880 4.180 4.180 ;
        RECT 3.880 2.540 4.180 4.180 ;
        RECT 2.160 2.540 4.180 2.840 ;
        RECT 2.330 3.880 2.630 4.820 ;
        RECT 2.190 4.480 2.590 6.480 ;
        RECT 2.160 0.840 2.460 2.850 ;
    END
  END S
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.840 -0.540 4.240 0.650 ;
        RECT 9.690 -0.540 11.590 0.650 ;
        RECT 15.840 -0.540 15.990 0.660 ;
        RECT 0.000 -0.540 17.160 0.540 ;
    END
  END GRND
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 4.690 7.270 8.090 8.460 ;
        RECT 0.000 7.380 17.160 8.460 ;
        RECT 13.710 7.270 16.110 8.460 ;
    END
  END POWR
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.080 3.260 15.380 6.290 ;
        RECT 15.770 1.900 16.170 2.700 ;
        RECT 15.080 3.260 16.120 3.560 ;
        RECT 15.820 1.900 16.120 3.560 ;
        RECT 15.080 4.090 15.720 4.490 ;
        RECT 14.780 5.090 15.380 6.290 ;
    END
  END CO
  OBS 
      LAYER Metal1 ;
        RECT 0.500 1.040 0.900 2.240 ;
        RECT 0.630 4.480 1.030 6.480 ;
        RECT 0.640 4.480 0.940 6.880 ;
        RECT 1.280 0.840 1.680 2.240 ;
        RECT 2.970 3.140 3.370 3.560 ;
        RECT 0.730 3.260 3.370 3.560 ;
        RECT 0.730 3.200 1.130 3.600 ;
        RECT 3.770 5.980 4.170 6.380 ;
        RECT 1.410 4.480 1.810 6.480 ;
        RECT 1.460 4.480 1.760 7.070 ;
        RECT 3.770 5.980 4.070 7.080 ;
        RECT 1.610 6.780 4.070 7.080 ;
        RECT 2.840 1.890 5.090 2.190 ;
        RECT 2.840 0.840 3.240 2.240 ;
        RECT 4.590 1.890 5.090 2.300 ;
        RECT 4.790 1.890 5.090 2.700 ;
        RECT 4.820 2.400 5.120 3.760 ;
        RECT 4.620 3.460 4.920 5.680 ;
        RECT 2.970 5.380 4.920 5.680 ;
        RECT 2.970 4.480 3.370 6.480 ;
        RECT 5.390 1.300 5.790 2.100 ;
        RECT 5.460 1.300 5.760 2.710 ;
        RECT 5.460 2.410 6.100 2.710 ;
        RECT 5.750 3.160 6.150 3.560 ;
        RECT 5.800 2.410 6.100 4.390 ;
        RECT 5.320 4.090 6.100 4.390 ;
        RECT 5.320 4.090 5.620 5.690 ;
        RECT 5.220 4.690 5.620 5.690 ;
        RECT 6.000 4.690 6.400 5.690 ;
        RECT 6.100 4.690 6.400 6.770 ;
        RECT 6.200 1.040 6.500 2.100 ;
        RECT 6.170 1.300 6.570 2.100 ;
        RECT 6.870 1.140 7.370 1.680 ;
        RECT 6.870 1.380 8.180 1.680 ;
        RECT 7.780 0.850 8.180 2.250 ;
        RECT 6.870 1.140 7.170 4.630 ;
        RECT 6.870 4.330 8.010 4.630 ;
        RECT 7.610 4.190 8.010 6.190 ;
        RECT 8.390 4.190 8.790 6.190 ;
        RECT 8.440 4.190 8.740 6.770 ;
        RECT 8.590 4.190 8.740 6.880 ;
        RECT 8.560 1.040 8.960 2.250 ;
        RECT 9.920 2.190 10.360 2.690 ;
        RECT 8.970 3.390 9.370 3.790 ;
        RECT 8.980 3.580 10.220 3.880 ;
        RECT 9.920 2.190 10.220 6.210 ;
        RECT 9.840 5.210 10.240 6.210 ;
        RECT 10.620 5.210 11.020 6.210 ;
        RECT 10.690 5.210 10.990 6.880 ;
        RECT 10.800 1.150 11.100 2.690 ;
        RECT 10.740 2.190 11.140 2.690 ;
        RECT 11.620 4.560 12.020 5.060 ;
        RECT 11.620 6.260 12.020 6.760 ;
        RECT 11.680 4.560 11.980 6.880 ;
        RECT 12.760 0.930 13.160 1.490 ;
        RECT 11.820 1.190 13.160 1.490 ;
        RECT 11.820 1.190 12.120 2.530 ;
        RECT 11.740 2.030 12.140 2.530 ;
        RECT 13.540 1.040 13.940 1.430 ;
        RECT 14.000 5.090 14.400 6.290 ;
        RECT 14.030 5.090 14.330 6.770 ;
        RECT 12.520 2.030 12.920 2.530 ;
        RECT 12.520 3.850 14.610 4.150 ;
        RECT 14.360 3.860 14.760 4.260 ;
        RECT 12.400 4.560 12.820 5.060 ;
        RECT 12.520 2.030 12.820 6.490 ;
        RECT 12.400 6.260 12.800 6.760 ;
        RECT 15.040 1.040 15.340 2.700 ;
        RECT 14.990 1.900 15.390 2.700 ;
  END 
END ADDHX1

MACRO CLKBUFX2
  CLASS  CORE ;
  FOREIGN CLKBUFX2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.960 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.120 2.770 1.800 3.170 ;
    END
  END A
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 -0.540 0.800 0.650 ;
        RECT 0.000 -0.540 3.960 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.330 0.900 2.630 6.670 ;
        RECT 2.330 3.430 3.120 3.830 ;
        RECT 2.280 5.170 2.680 6.670 ;
        RECT 2.280 0.900 2.680 2.250 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 7.380 3.960 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 1.300 5.170 1.900 6.670 ;
        RECT 1.300 4.680 1.700 6.880 ;
        RECT 1.300 1.040 1.900 2.250 ;
        RECT 0.520 1.250 0.920 2.250 ;
        RECT 0.520 3.920 2.030 4.220 ;
        RECT 1.630 3.880 2.030 4.280 ;
        RECT 0.520 1.250 0.820 7.080 ;
        RECT 0.520 4.680 0.920 7.080 ;
        RECT 3.060 5.170 3.460 6.880 ;
  END 
END CLKBUFX2

MACRO CLKBUFX3
  CLASS  CORE ;
  FOREIGN CLKBUFX3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.960 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.840 2.810 1.460 3.210 ;
    END
  END A
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 -0.540 3.440 0.650 ;
        RECT 0.000 -0.540 3.960 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.260 1.250 2.660 2.150 ;
        RECT 2.770 2.750 3.170 3.170 ;
        RECT 2.360 3.770 3.080 4.070 ;
        RECT 2.780 2.450 3.080 4.070 ;
        RECT 2.360 2.450 3.080 2.750 ;
        RECT 2.260 4.370 2.660 6.670 ;
        RECT 2.360 3.770 2.660 6.670 ;
        RECT 2.360 1.250 2.660 2.750 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 7.380 3.960 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 1.280 4.280 1.680 6.880 ;
        RECT 1.280 4.370 1.880 6.880 ;
        RECT 1.280 1.150 1.880 2.150 ;
        RECT 1.280 1.150 1.680 2.410 ;
        RECT 0.500 1.250 0.900 2.410 ;
        RECT 0.190 2.110 0.900 2.410 ;
        RECT 1.760 3.060 2.360 3.460 ;
        RECT 0.190 2.110 0.490 3.980 ;
        RECT 1.760 3.060 2.060 3.980 ;
        RECT 0.190 3.680 2.060 3.980 ;
        RECT 0.500 3.680 0.800 7.080 ;
        RECT 0.500 4.280 0.900 7.080 ;
        RECT 3.040 4.370 3.440 6.880 ;
        RECT 3.040 1.150 3.440 2.150 ;
  END 
END CLKBUFX3

MACRO CLKBUFX1
  CLASS  CORE ;
  FOREIGN CLKBUFX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.300 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.790 3.430 1.190 4.090 ;
        RECT 0.790 3.690 1.500 4.090 ;
    END
  END A
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 -0.540 2.500 0.650 ;
        RECT 0.000 -0.540 3.300 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.260 1.250 2.660 2.050 ;
        RECT 2.260 4.490 2.660 6.670 ;
        RECT 2.360 1.250 2.660 6.670 ;
        RECT 2.110 3.430 2.660 3.830 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 7.270 2.500 8.460 ;
        RECT 0.000 7.380 3.300 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 1.480 4.490 1.880 6.770 ;
        RECT 1.280 4.850 1.880 6.770 ;
        RECT 1.280 1.150 1.880 1.900 ;
        RECT 1.480 1.150 1.880 2.050 ;
        RECT 0.500 1.250 0.900 1.900 ;
        RECT 0.500 1.250 0.800 2.750 ;
        RECT 0.190 2.450 2.060 2.750 ;
        RECT 1.660 2.450 2.060 2.850 ;
        RECT 0.190 2.450 0.490 5.150 ;
        RECT 0.190 4.850 0.900 5.150 ;
        RECT 0.500 4.850 0.900 6.670 ;
  END 
END CLKBUFX1

MACRO DFFSRX1
  CLASS  CORE ;
  FOREIGN DFFSRX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.460 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 17.770 1.730 18.170 2.380 ;
        RECT 17.870 2.770 18.350 3.170 ;
        RECT 17.770 4.850 18.170 6.670 ;
        RECT 17.870 1.730 18.170 6.670 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 19.320 3.480 19.680 3.780 ;
        RECT 19.330 4.850 19.730 6.670 ;
        RECT 19.330 1.730 19.730 2.380 ;
        RECT 19.380 1.730 19.680 6.670 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.680 1.250 0.980 6.190 ;
        RECT 0.680 2.770 1.190 3.170 ;
        RECT 0.630 4.370 1.030 6.190 ;
        RECT 0.630 1.250 1.030 1.900 ;
    END
  END D
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 -0.540 3.700 0.650 ;
        RECT 0.000 -0.540 20.460 0.540 ;
        RECT 15.770 -0.540 19.960 0.650 ;
    END
  END GRND
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.070 0.840 7.470 1.240 ;
        RECT 15.070 0.840 15.470 1.240 ;
        RECT 7.070 0.840 15.470 1.140 ;
        RECT 8.050 0.840 8.450 1.850 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.290 2.770 5.150 3.170 ;
    END
  END CK
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 7.270 2.100 8.460 ;
        RECT 0.000 7.380 20.460 8.460 ;
        RECT 18.600 7.270 19.950 8.460 ;
        RECT 10.070 7.270 13.270 8.460 ;
    END
  END POWR
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.810 6.580 8.210 7.080 ;
        RECT 14.330 6.580 14.730 7.080 ;
        RECT 7.810 6.580 14.730 6.880 ;
        RECT 8.710 6.070 9.110 6.880 ;
    END
  END SN
  OBS 
      LAYER Metal1 ;
        RECT 1.410 1.250 1.810 1.900 ;
        RECT 1.410 4.370 1.810 6.190 ;
        RECT 1.510 1.250 1.810 6.970 ;
        RECT 1.510 6.670 3.690 6.970 ;
        RECT 3.290 6.670 3.690 7.080 ;
        RECT 3.590 1.250 3.990 1.900 ;
        RECT 2.990 3.660 3.390 4.060 ;
        RECT 2.990 3.760 3.990 4.060 ;
        RECT 3.690 1.250 3.990 4.860 ;
        RECT 3.590 4.460 3.990 4.860 ;
        RECT 4.370 5.880 4.770 6.280 ;
        RECT 4.420 5.880 4.720 6.880 ;
        RECT 4.410 1.040 4.710 1.900 ;
        RECT 4.370 1.250 4.770 1.900 ;
        RECT 6.470 1.040 6.770 2.090 ;
        RECT 6.470 1.790 7.730 2.090 ;
        RECT 7.330 1.790 7.730 2.440 ;
        RECT 5.770 1.790 6.170 2.440 ;
        RECT 5.770 2.740 8.810 3.040 ;
        RECT 8.410 2.740 8.810 3.240 ;
        RECT 5.770 1.790 6.070 4.760 ;
        RECT 5.770 4.460 6.950 4.760 ;
        RECT 6.550 4.460 6.950 4.860 ;
        RECT 8.060 5.160 9.290 5.460 ;
        RECT 8.890 5.160 9.290 5.560 ;
        RECT 8.060 5.160 8.360 6.180 ;
        RECT 5.770 5.880 8.360 6.180 ;
        RECT 5.770 5.880 7.730 6.280 ;
        RECT 7.110 5.880 7.510 6.880 ;
        RECT 2.190 1.250 2.590 1.900 ;
        RECT 8.890 1.790 9.290 2.440 ;
        RECT 2.190 1.250 2.490 6.190 ;
        RECT 9.110 2.140 9.410 4.760 ;
        RECT 7.250 4.460 9.410 4.760 ;
        RECT 8.110 4.460 8.510 4.860 ;
        RECT 7.250 4.460 7.550 5.460 ;
        RECT 2.190 5.160 7.550 5.460 ;
        RECT 2.190 4.370 2.590 6.190 ;
        RECT 10.290 1.500 10.690 1.910 ;
        RECT 9.890 2.840 10.590 3.240 ;
        RECT 10.290 1.500 10.590 6.190 ;
        RECT 10.290 4.370 10.690 6.190 ;
        RECT 11.070 1.500 11.470 1.910 ;
        RECT 11.080 3.570 12.550 3.870 ;
        RECT 12.150 3.570 12.550 3.970 ;
        RECT 11.080 1.500 11.380 6.190 ;
        RECT 11.070 4.370 11.470 6.190 ;
        RECT 15.770 1.150 16.070 2.090 ;
        RECT 14.810 1.790 16.070 2.090 ;
        RECT 14.810 1.790 15.210 2.440 ;
        RECT 13.250 1.790 13.650 2.440 ;
        RECT 13.250 2.140 14.330 2.440 ;
        RECT 14.030 2.740 16.290 3.040 ;
        RECT 15.890 2.740 16.290 3.240 ;
        RECT 14.030 2.140 14.330 4.860 ;
        RECT 14.030 4.460 14.430 4.860 ;
        RECT 13.250 5.880 16.770 6.280 ;
        RECT 15.030 5.880 15.430 6.880 ;
        RECT 11.850 1.500 12.250 1.910 ;
        RECT 16.370 1.790 16.770 2.440 ;
        RECT 11.950 1.500 12.250 3.270 ;
        RECT 11.950 2.970 13.150 3.270 ;
        RECT 12.850 2.970 13.150 4.670 ;
        RECT 11.850 4.370 13.150 4.670 ;
        RECT 16.590 2.140 16.890 4.760 ;
        RECT 15.590 4.460 16.890 4.760 ;
        RECT 15.590 4.460 15.990 5.580 ;
        RECT 11.850 5.280 15.990 5.580 ;
        RECT 11.850 4.370 12.250 6.190 ;
        RECT 18.550 4.850 18.950 6.670 ;
        RECT 18.600 4.850 18.900 6.770 ;
        RECT 18.600 1.150 18.900 2.380 ;
        RECT 18.550 1.730 18.950 2.380 ;
  END 
END DFFSRX1

MACRO DFFX1
  CLASS  CORE ;
  FOREIGN DFFX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.480 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 15.210 1.420 15.510 6.670 ;
        RECT 16.020 3.270 16.640 3.670 ;
        RECT 16.020 2.770 16.320 3.670 ;
        RECT 15.210 2.770 16.320 3.070 ;
        RECT 15.160 4.070 15.560 6.670 ;
        RECT 15.160 1.420 15.560 2.420 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.720 1.420 17.120 2.420 ;
        RECT 16.940 2.820 17.640 3.120 ;
        RECT 16.940 2.120 17.240 4.370 ;
        RECT 16.720 4.070 17.120 6.670 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.760 3.430 2.460 3.830 ;
    END
  END D
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.270 -0.540 17.480 0.650 ;
        RECT 0.000 -0.540 18.480 0.540 ;
    END
  END GRND
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.780 2.820 1.180 3.520 ;
    END
  END CK
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.940 7.270 17.150 8.460 ;
        RECT 0.000 7.380 18.480 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.260 0.840 0.850 1.240 ;
        RECT 0.550 0.840 0.850 2.330 ;
        RECT 0.550 1.730 0.950 2.330 ;
        RECT 0.180 2.030 0.950 2.330 ;
        RECT 0.180 2.030 0.480 4.790 ;
        RECT 0.180 4.490 0.950 4.790 ;
        RECT 0.550 4.490 0.950 6.190 ;
        RECT 1.330 4.490 1.730 6.770 ;
        RECT 1.330 1.150 1.730 2.330 ;
        RECT 2.110 1.730 2.510 2.330 ;
        RECT 3.510 1.730 3.910 2.330 ;
        RECT 2.110 2.030 3.910 2.330 ;
        RECT 2.860 2.030 3.160 4.790 ;
        RECT 2.110 4.490 3.910 4.790 ;
        RECT 2.110 4.490 2.510 6.190 ;
        RECT 3.510 4.490 3.910 6.190 ;
        RECT 4.290 1.730 4.690 2.330 ;
        RECT 4.390 3.760 5.770 4.060 ;
        RECT 5.370 3.690 5.770 4.090 ;
        RECT 4.390 1.730 4.690 6.190 ;
        RECT 4.290 4.490 4.690 6.190 ;
        RECT 7.460 5.790 7.860 6.770 ;
        RECT 7.460 1.150 7.860 2.330 ;
        RECT 6.680 1.730 7.080 2.330 ;
        RECT 6.780 3.260 8.040 3.560 ;
        RECT 7.640 3.210 8.040 3.610 ;
        RECT 6.780 1.730 7.080 4.890 ;
        RECT 6.680 4.490 7.080 4.890 ;
        RECT 5.070 1.730 5.470 2.330 ;
        RECT 8.240 1.730 8.640 2.330 ;
        RECT 5.070 2.030 6.380 2.330 ;
        RECT 9.640 1.730 10.040 2.330 ;
        RECT 8.240 2.030 10.040 2.330 ;
        RECT 8.240 4.490 10.040 4.790 ;
        RECT 6.080 2.030 6.380 5.490 ;
        RECT 5.070 5.190 8.640 5.490 ;
        RECT 5.070 4.490 5.470 6.190 ;
        RECT 8.340 1.730 8.640 6.190 ;
        RECT 8.240 4.490 8.640 6.190 ;
        RECT 9.640 4.490 10.040 6.190 ;
        RECT 10.420 1.730 10.820 2.330 ;
        RECT 10.520 3.070 11.700 3.370 ;
        RECT 11.300 3.020 11.700 3.420 ;
        RECT 10.520 1.730 10.820 6.190 ;
        RECT 10.420 4.490 10.820 6.190 ;
        RECT 13.380 5.790 13.780 6.770 ;
        RECT 13.380 1.150 13.780 2.330 ;
        RECT 12.600 1.730 13.000 2.330 ;
        RECT 12.700 3.250 13.960 3.550 ;
        RECT 13.560 3.210 13.960 3.610 ;
        RECT 12.700 1.730 13.000 4.890 ;
        RECT 12.600 4.490 13.000 4.890 ;
        RECT 11.200 1.730 11.600 2.330 ;
        RECT 11.200 2.030 12.300 2.330 ;
        RECT 14.160 1.730 14.560 2.330 ;
        RECT 14.260 2.820 14.860 3.220 ;
        RECT 12.000 2.030 12.300 5.490 ;
        RECT 11.200 5.190 14.560 5.490 ;
        RECT 11.200 4.490 11.600 6.190 ;
        RECT 14.260 1.730 14.560 6.190 ;
        RECT 14.160 4.490 14.560 6.190 ;
        RECT 15.940 4.070 16.340 6.770 ;
        RECT 15.940 1.150 16.340 2.420 ;
  END 
END DFFX1

MACRO MX2X1
  CLASS  CORE ;
  FOREIGN MX2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.920 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.620 2.830 6.020 3.230 ;
        RECT 5.960 2.770 6.420 3.170 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.840 2.160 1.140 2.710 ;
        RECT 1.460 2.410 1.860 2.810 ;
        RECT 0.790 2.410 1.860 2.710 ;
    END
  END B
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 4.620 -0.540 5.020 0.660 ;
        RECT 6.700 -0.540 6.980 0.660 ;
        RECT 0.000 -0.540 7.920 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.680 3.580 6.980 6.270 ;
        RECT 6.780 2.220 7.080 3.880 ;
        RECT 6.580 4.450 6.980 6.270 ;
        RECT 6.580 1.260 6.980 1.910 ;
        RECT 6.640 1.260 6.940 2.520 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.840 7.270 4.240 8.460 ;
        RECT 6.780 7.270 7.180 8.460 ;
        RECT 0.000 7.380 7.920 8.460 ;
    END
  END POWR
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.980 4.050 1.380 4.450 ;
        RECT 1.010 4.090 1.800 4.490 ;
    END
  END S0
  OBS 
      LAYER Metal1 ;
        RECT 1.280 4.850 1.680 6.880 ;
        RECT 1.280 1.040 1.680 1.590 ;
        RECT 0.500 0.940 0.900 1.590 ;
        RECT 0.150 1.290 0.900 1.590 ;
        RECT 0.150 3.120 2.760 3.420 ;
        RECT 2.360 3.090 2.760 3.490 ;
        RECT 0.150 1.290 0.450 5.150 ;
        RECT 0.150 4.850 0.900 5.150 ;
        RECT 0.500 4.850 0.900 6.670 ;
        RECT 2.060 0.940 2.460 1.590 ;
        RECT 2.160 0.940 2.460 2.790 ;
        RECT 2.160 2.490 3.360 2.790 ;
        RECT 3.060 2.490 3.360 4.550 ;
        RECT 2.160 4.250 3.360 4.550 ;
        RECT 2.160 4.250 2.460 6.670 ;
        RECT 2.060 4.850 2.460 6.670 ;
        RECT 2.840 0.940 3.240 1.590 ;
        RECT 2.940 0.940 3.240 2.190 ;
        RECT 2.940 1.890 3.960 2.190 ;
        RECT 3.660 1.890 3.960 5.150 ;
        RECT 2.840 4.850 3.960 5.150 ;
        RECT 2.840 4.850 3.240 6.670 ;
        RECT 2.840 6.370 4.120 6.670 ;
        RECT 3.820 6.670 5.110 6.970 ;
        RECT 4.710 6.670 5.110 7.070 ;
        RECT 3.620 0.940 4.020 1.590 ;
        RECT 3.620 1.290 5.420 1.590 ;
        RECT 5.020 1.260 5.420 1.910 ;
        RECT 5.020 1.260 5.320 6.270 ;
        RECT 3.620 5.450 5.420 5.750 ;
        RECT 3.620 5.450 4.020 5.850 ;
        RECT 5.020 4.450 5.420 6.270 ;
        RECT 5.800 4.450 6.200 6.880 ;
        RECT 5.800 1.040 6.200 1.910 ;
  END 
END MX2X1

MACRO XOR2X1
  CLASS  CORE ;
  FOREIGN XOR2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.260 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.090 3.430 4.490 3.880 ;
        RECT 4.090 3.480 5.120 3.880 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.980 2.530 1.380 3.130 ;
        RECT 5.620 3.480 6.020 3.880 ;
        RECT 5.620 2.830 5.920 3.880 ;
        RECT 5.390 2.770 5.810 3.150 ;
        RECT 0.980 2.830 5.920 3.130 ;
    END
  END B
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.540 7.260 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.240 1.250 4.640 2.090 ;
        RECT 5.020 4.280 6.620 4.580 ;
        RECT 6.320 1.790 6.620 4.580 ;
        RECT 6.070 1.790 6.620 2.510 ;
        RECT 4.240 1.790 6.620 2.090 ;
        RECT 5.020 4.280 5.420 6.280 ;
        RECT 4.440 0.840 4.840 1.490 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.840 7.270 2.840 8.460 ;
        RECT 0.000 7.380 7.260 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 1.280 4.070 1.680 6.670 ;
        RECT 1.280 1.040 1.680 1.490 ;
        RECT 2.060 4.070 2.460 6.770 ;
        RECT 0.500 0.840 0.900 2.090 ;
        RECT 2.060 0.840 2.460 2.090 ;
        RECT 0.380 1.790 3.060 2.090 ;
        RECT 2.660 1.790 3.060 2.290 ;
        RECT 0.380 1.790 0.680 3.770 ;
        RECT 0.380 3.470 3.790 3.770 ;
        RECT 3.390 3.470 3.790 3.880 ;
        RECT 0.500 3.470 0.900 6.670 ;
        RECT 3.460 4.280 3.860 6.880 ;
        RECT 3.460 1.040 3.860 1.900 ;
        RECT 5.220 0.840 5.620 1.490 ;
        RECT 4.240 4.280 4.640 7.080 ;
        RECT 5.800 5.080 6.200 7.080 ;
        RECT 4.240 6.680 6.200 7.080 ;
        RECT 6.000 1.040 6.400 1.490 ;
  END 
END XOR2X1

MACRO OAI33X1
  CLASS  CORE ;
  FOREIGN OAI33X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.560 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.090 2.820 4.490 3.400 ;
        RECT 3.740 3.000 4.490 3.400 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.410 2.990 5.810 3.780 ;
    END
  END A1
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 7.520 -0.540 9.920 0.650 ;
        RECT 0.000 -0.540 10.560 0.540 ;
    END
  END GRND
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.340 3.430 6.740 4.080 ;
        RECT 6.340 3.430 7.080 3.830 ;
    END
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 9.660 1.250 10.060 2.350 ;
        RECT 9.660 4.250 10.060 7.080 ;
        RECT 9.760 1.250 10.060 7.080 ;
        RECT 9.370 3.430 10.060 3.830 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.700 3.200 3.170 3.600 ;
        RECT 2.770 3.200 3.170 3.780 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.760 3.200 2.160 3.830 ;
        RECT 1.450 3.430 2.160 3.830 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.380 2.490 0.780 3.170 ;
        RECT 0.380 2.770 1.190 3.170 ;
    END
  END B2
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 6.880 7.270 7.680 8.460 ;
        RECT 0.000 7.380 10.560 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.500 4.480 1.500 6.880 ;
        RECT 0.500 1.040 1.500 2.090 ;
        RECT 1.880 4.480 2.280 7.080 ;
        RECT 2.660 4.480 3.060 7.080 ;
        RECT 2.660 1.040 3.060 2.090 ;
        RECT 4.220 4.480 4.620 7.080 ;
        RECT 5.000 4.480 5.400 7.080 ;
        RECT 4.060 0.840 5.920 1.140 ;
        RECT 1.880 1.440 2.280 2.090 ;
        RECT 4.060 0.840 4.360 2.090 ;
        RECT 3.440 1.440 4.360 2.090 ;
        RECT 5.620 0.840 5.920 2.090 ;
        RECT 5.520 1.440 5.920 2.090 ;
        RECT 1.980 1.440 2.280 2.700 ;
        RECT 3.440 1.440 3.740 2.700 ;
        RECT 1.980 2.400 3.740 2.700 ;
        RECT 5.780 4.480 6.180 6.880 ;
        RECT 4.740 1.440 5.140 2.090 ;
        RECT 6.300 1.440 6.700 2.090 ;
        RECT 6.300 1.440 6.600 2.690 ;
        RECT 4.790 2.390 7.300 2.690 ;
        RECT 6.900 2.390 7.300 2.890 ;
        RECT 4.790 1.440 5.090 4.180 ;
        RECT 3.540 3.880 5.090 4.180 ;
        RECT 3.540 3.880 3.840 7.080 ;
        RECT 3.440 4.480 3.840 7.080 ;
        RECT 7.700 1.700 8.100 2.350 ;
        RECT 7.800 2.750 9.180 3.050 ;
        RECT 8.780 2.750 9.180 3.150 ;
        RECT 7.800 1.700 8.100 6.670 ;
        RECT 7.700 4.850 8.100 6.670 ;
        RECT 8.880 4.250 9.280 6.880 ;
        RECT 8.480 4.850 9.280 6.880 ;
        RECT 8.480 1.150 9.280 2.350 ;
  END 
END OAI33X1

MACRO OAI22X1
  CLASS  CORE ;
  FOREIGN OAI22X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.920 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.480 3.640 2.880 4.490 ;
        RECT 2.110 4.090 2.880 4.490 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.430 3.430 3.830 4.450 ;
        RECT 3.430 4.050 3.840 4.450 ;
    END
  END A1
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 -0.540 1.680 0.650 ;
        RECT 0.000 -0.540 7.920 0.540 ;
        RECT 4.750 -0.540 7.150 0.650 ;
        RECT 0.500 -0.540 1.700 0.640 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.780 1.250 7.180 2.350 ;
        RECT 6.780 4.250 7.180 7.080 ;
        RECT 6.880 1.250 7.180 7.080 ;
        RECT 6.730 2.770 7.180 3.170 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 2.990 1.850 3.830 ;
        RECT 1.450 2.990 1.980 3.390 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.680 4.050 1.080 4.450 ;
        RECT 0.780 4.090 1.180 4.490 ;
    END
  END B1
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 7.270 4.040 8.460 ;
        RECT 0.000 7.380 7.920 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.500 4.850 0.900 6.770 ;
        RECT 1.280 4.850 1.680 6.670 ;
        RECT 1.280 1.150 1.680 2.090 ;
        RECT 2.840 5.800 3.240 6.670 ;
        RECT 3.620 5.800 4.020 6.770 ;
        RECT 2.160 0.840 3.920 1.140 ;
        RECT 3.620 0.840 3.920 2.090 ;
        RECT 0.500 1.440 0.900 2.090 ;
        RECT 2.160 0.840 2.460 2.090 ;
        RECT 3.620 1.440 4.020 2.090 ;
        RECT 0.600 1.440 0.900 2.690 ;
        RECT 2.060 1.440 2.360 2.690 ;
        RECT 0.600 2.390 2.360 2.690 ;
        RECT 2.840 1.440 3.240 2.090 ;
        RECT 2.940 1.440 3.240 2.690 ;
        RECT 2.940 2.390 4.820 2.690 ;
        RECT 4.420 2.390 4.820 3.090 ;
        RECT 4.420 2.390 4.720 5.150 ;
        RECT 2.060 4.850 4.720 5.150 ;
        RECT 2.060 4.850 2.460 6.670 ;
        RECT 6.000 4.250 6.400 6.880 ;
        RECT 5.800 5.260 6.400 6.880 ;
        RECT 5.800 1.150 6.400 1.900 ;
        RECT 6.000 1.150 6.400 2.350 ;
        RECT 5.020 1.250 5.420 1.900 ;
        RECT 6.100 3.450 6.500 3.850 ;
        RECT 5.120 3.550 6.500 3.850 ;
        RECT 5.120 1.250 5.420 7.080 ;
        RECT 5.020 5.260 5.420 7.080 ;
  END 
END OAI22X1

MACRO OAI21X1
  CLASS  CORE ;
  FOREIGN OAI21X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.850 2.700 2.250 3.170 ;
        RECT 1.850 2.770 2.460 3.170 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.740 2.770 1.140 3.580 ;
    END
  END A1
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 4.010 -0.540 4.410 0.650 ;
        RECT 0.000 -0.540 5.280 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.020 0.840 3.320 7.080 ;
        RECT 3.020 2.110 3.830 2.510 ;
        RECT 3.010 0.840 3.410 1.580 ;
        RECT 2.930 3.980 3.330 7.080 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.090 2.770 4.490 3.580 ;
        RECT 3.620 3.180 4.490 3.580 ;
    END
  END B0
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.670 3.980 1.770 8.460 ;
        RECT 0.000 7.380 5.280 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 1.450 1.040 1.850 1.580 ;
        RECT 2.150 3.980 2.550 7.080 ;
        RECT 0.670 0.840 1.070 1.580 ;
        RECT 2.230 0.840 2.630 1.580 ;
        RECT 0.770 0.840 1.070 2.180 ;
        RECT 2.230 0.840 2.530 2.180 ;
        RECT 0.770 1.880 2.530 2.180 ;
        RECT 3.710 3.980 4.110 6.880 ;
  END 
END OAI21X1

MACRO AOI22X1
  CLASS  CORE ;
  FOREIGN AOI22X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 1.940 1.850 2.510 ;
        RECT 1.450 1.940 2.100 2.340 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 2.770 1.190 3.170 ;
    END
  END A1
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.540 5.280 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.520 3.670 1.920 5.350 ;
        RECT 1.620 3.070 2.700 3.370 ;
        RECT 2.400 0.840 2.700 3.370 ;
        RECT 2.160 2.820 2.700 3.370 ;
        RECT 2.300 0.840 2.700 1.540 ;
        RECT 1.300 4.080 1.920 5.350 ;
        RECT 1.620 3.070 1.920 5.350 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.000 2.770 3.400 3.170 ;
        RECT 3.430 3.430 3.830 3.830 ;
        RECT 3.430 2.870 3.730 3.830 ;
        RECT 3.000 2.870 3.730 3.170 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.090 2.770 4.630 3.170 ;
    END
  END B1
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.300 7.270 2.580 8.460 ;
        RECT 0.000 7.380 5.280 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.520 1.040 0.920 1.540 ;
        RECT 1.300 0.840 1.920 1.540 ;
        RECT 3.080 4.950 3.880 6.880 ;
        RECT 3.080 0.840 3.480 1.540 ;
        RECT 3.480 1.240 3.880 1.950 ;
        RECT 2.300 4.130 4.660 4.530 ;
        RECT 2.300 3.670 2.700 6.670 ;
        RECT 0.520 6.270 2.700 6.670 ;
        RECT 0.520 4.080 0.920 7.080 ;
        RECT 4.260 4.080 4.660 7.080 ;
        RECT 4.260 1.040 4.660 1.950 ;
  END 
END AOI22X1

MACRO AOI21X1
  CLASS  CORE ;
  FOREIGN AOI21X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.960 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.580 3.270 1.980 3.830 ;
        RECT 1.580 3.430 2.510 3.830 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.680 2.350 1.080 3.830 ;
        RECT 0.680 3.430 1.190 3.830 ;
    END
  END A1
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.540 3.960 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.060 1.250 2.460 1.950 ;
        RECT 2.840 4.070 3.240 6.670 ;
        RECT 2.840 2.710 3.140 6.670 ;
        RECT 2.820 2.710 3.140 3.120 ;
        RECT 2.160 2.710 3.140 3.010 ;
        RECT 2.260 0.840 2.660 1.540 ;
        RECT 2.160 1.250 2.460 3.010 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.860 1.940 3.260 2.390 ;
        RECT 3.480 2.090 3.780 2.460 ;
        RECT 2.860 2.090 3.780 2.390 ;
    END
  END B0
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 7.270 3.300 8.460 ;
        RECT 0.000 7.380 3.960 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.500 1.040 0.900 1.950 ;
        RECT 1.280 4.950 1.680 6.770 ;
        RECT 1.280 1.250 1.680 1.950 ;
        RECT 0.500 4.250 2.460 4.650 ;
        RECT 0.500 4.250 0.900 6.670 ;
        RECT 2.060 4.250 2.460 6.670 ;
        RECT 3.040 1.040 3.440 1.540 ;
  END 
END AOI21X1

MACRO FILL4
  CLASS  CORE ;
  FOREIGN FILL4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.640 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.120 -0.540 1.520 0.650 ;
        RECT 0.000 -0.540 2.640 0.540 ;
    END
  END GRND
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.020 7.170 1.620 8.460 ;
        RECT 0.000 7.380 2.640 8.460 ;
    END
  END POWR
END FILL4

MACRO FILL2
  CLASS  CORE ;
  FOREIGN FILL2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.320 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.540 1.320 0.540 ;
    END
  END GRND
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 7.380 1.320 8.460 ;
    END
  END POWR
END FILL2

MACRO FILL1
  CLASS  CORE ;
  FOREIGN FILL1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.660 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.540 0.660 0.540 ;
    END
  END GRND
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 7.380 0.660 8.460 ;
    END
  END POWR
END FILL1

MACRO BUFX3
  CLASS  CORE ;
  FOREIGN BUFX3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.960 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.150 2.390 1.800 2.790 ;
        RECT 1.500 2.390 1.800 3.120 ;
    END
  END A
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 -0.540 0.800 0.650 ;
        RECT 0.000 -0.540 3.960 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.340 0.840 2.640 7.080 ;
        RECT 2.340 2.770 3.120 3.170 ;
        RECT 2.280 4.280 2.680 7.080 ;
        RECT 2.280 0.840 2.680 1.990 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 7.270 0.800 8.460 ;
        RECT 0.000 7.380 3.960 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 1.500 4.280 1.900 6.880 ;
        RECT 1.300 4.870 1.900 6.880 ;
        RECT 1.300 1.040 1.900 1.990 ;
        RECT 0.520 1.290 0.920 1.990 ;
        RECT 1.640 3.480 2.040 3.880 ;
        RECT 0.550 3.580 2.040 3.880 ;
        RECT 0.550 1.290 0.850 6.670 ;
        RECT 0.520 4.870 0.920 6.670 ;
        RECT 3.060 4.280 3.460 6.880 ;
        RECT 3.060 1.040 3.460 1.990 ;
  END 
END BUFX3

MACRO OR4X1
  CLASS  CORE ;
  FOREIGN OR4X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.240 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.680 3.860 1.080 4.260 ;
        RECT 0.770 3.430 1.190 3.860 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 2.390 1.850 3.170 ;
        RECT 1.450 2.390 2.000 2.790 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.750 2.390 5.150 3.170 ;
        RECT 4.750 2.390 5.160 2.790 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.070 3.430 6.470 4.260 ;
        RECT 6.070 3.860 6.540 4.260 ;
    END
  END D
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.070 -0.540 3.470 0.650 ;
        RECT 6.840 -0.540 8.440 0.650 ;
        RECT 0.000 -0.540 9.240 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 8.020 1.250 8.420 6.670 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 7.260 1.820 8.460 ;
        RECT 0.000 7.380 9.240 8.460 ;
        RECT 4.960 7.270 8.560 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.500 1.040 0.900 1.490 ;
        RECT 1.420 5.460 1.820 6.760 ;
        RECT 2.060 1.040 2.460 1.490 ;
        RECT 0.640 4.660 2.800 5.060 ;
        RECT 0.640 4.660 1.040 6.660 ;
        RECT 2.200 4.660 2.800 6.660 ;
        RECT 2.400 2.870 2.800 7.070 ;
        RECT 3.180 2.870 3.580 7.070 ;
        RECT 4.280 1.040 4.680 1.490 ;
        RECT 3.960 4.660 4.560 6.660 ;
        RECT 5.720 4.660 6.120 6.660 ;
        RECT 3.960 6.260 6.120 6.660 ;
        RECT 3.960 2.870 4.360 7.070 ;
        RECT 5.840 1.040 6.240 1.490 ;
        RECT 7.240 4.490 7.640 6.770 ;
        RECT 7.240 1.150 7.640 2.050 ;
        RECT 1.280 0.840 1.680 1.490 ;
        RECT 5.060 0.840 5.460 1.490 ;
        RECT 1.380 0.840 1.680 2.090 ;
        RECT 5.100 0.840 5.400 2.090 ;
        RECT 1.380 1.790 5.760 2.090 ;
        RECT 5.460 2.450 7.710 2.750 ;
        RECT 7.310 2.450 7.710 2.850 ;
        RECT 5.460 1.790 5.760 4.360 ;
        RECT 5.030 4.060 5.760 4.360 ;
        RECT 5.030 4.060 5.330 5.860 ;
        RECT 4.940 4.660 5.340 5.860 ;
  END 
END OR4X1

MACRO OR2X1
  CLASS  CORE ;
  FOREIGN OR2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.960 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 4.090 2.090 4.490 ;
        RECT 2.090 3.550 2.490 3.950 ;
        RECT 2.090 3.550 2.390 4.440 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 2.300 1.100 3.170 ;
        RECT 0.700 2.770 1.190 3.170 ;
    END
  END B
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.600 -0.540 3.430 0.650 ;
        RECT 0.000 -0.540 3.960 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.940 1.250 3.340 1.900 ;
        RECT 3.180 1.600 3.480 5.150 ;
        RECT 2.940 4.850 3.340 6.670 ;
        RECT 2.770 4.090 3.480 4.490 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.630 7.270 3.430 8.460 ;
        RECT 0.000 7.380 3.960 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.600 1.150 1.000 1.900 ;
        RECT 1.380 4.850 1.780 6.670 ;
        RECT 2.160 4.850 2.560 6.770 ;
        RECT 2.160 1.150 2.560 1.900 ;
        RECT 1.380 1.250 1.780 1.900 ;
        RECT 1.480 1.250 1.780 2.500 ;
        RECT 1.490 2.200 2.860 2.630 ;
        RECT 2.460 2.200 2.860 2.700 ;
        RECT 1.490 2.200 1.790 3.770 ;
        RECT 0.600 3.470 1.790 3.770 ;
        RECT 0.600 3.470 0.900 6.670 ;
        RECT 0.600 4.850 1.000 6.670 ;
  END 
END OR2X1

MACRO NOR4X1
  CLASS  CORE ;
  FOREIGN NOR4X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.540 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.840 2.110 1.990 2.510 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.790 2.770 3.780 3.170 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.460 2.770 6.510 3.170 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 7.410 2.110 8.400 2.510 ;
    END
  END D
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 3.970 -0.540 5.170 0.650 ;
        RECT 8.490 -0.540 8.890 0.850 ;
        RECT 0.000 -0.540 12.540 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 11.430 0.840 11.830 1.920 ;
        RECT 11.430 4.260 11.830 7.080 ;
        RECT 11.530 0.840 11.830 7.080 ;
        RECT 11.400 3.480 11.830 3.780 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.730 7.270 1.930 8.460 ;
        RECT 4.430 7.270 4.830 8.460 ;
        RECT 8.960 7.270 9.760 8.460 ;
        RECT 0.000 7.380 12.540 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 1.410 4.280 1.810 6.770 ;
        RECT 1.410 1.040 1.810 1.490 ;
        RECT 2.970 1.040 3.370 1.490 ;
        RECT 0.730 3.680 2.490 3.980 ;
        RECT 0.730 3.680 1.030 6.480 ;
        RECT 0.630 4.280 1.030 6.480 ;
        RECT 2.190 3.680 2.490 6.480 ;
        RECT 3.750 4.280 4.150 6.480 ;
        RECT 2.290 4.280 2.590 7.080 ;
        RECT 3.750 4.280 4.050 7.080 ;
        RECT 2.290 6.780 4.050 7.080 ;
        RECT 3.070 3.680 6.230 3.980 ;
        RECT 5.930 3.680 6.230 6.480 ;
        RECT 3.070 3.680 3.370 6.480 ;
        RECT 2.970 4.280 3.370 6.480 ;
        RECT 5.930 4.280 6.330 6.480 ;
        RECT 5.930 1.040 6.330 1.490 ;
        RECT 7.490 1.040 7.890 1.490 ;
        RECT 5.150 4.280 5.550 6.480 ;
        RECT 6.710 4.280 7.110 6.480 ;
        RECT 8.270 4.280 8.670 6.480 ;
        RECT 5.170 4.280 5.470 7.080 ;
        RECT 6.780 4.280 7.080 7.080 ;
        RECT 8.360 4.280 8.660 7.080 ;
        RECT 5.170 6.780 8.660 7.080 ;
        RECT 2.190 0.840 2.590 1.490 ;
        RECT 6.710 0.840 7.110 1.490 ;
        RECT 2.290 0.840 2.590 2.090 ;
        RECT 2.290 1.790 7.110 2.090 ;
        RECT 6.810 0.840 7.110 3.840 ;
        RECT 6.810 3.540 9.420 3.840 ;
        RECT 9.020 3.480 9.420 3.880 ;
        RECT 7.540 3.540 7.840 6.480 ;
        RECT 7.490 4.280 7.890 6.480 ;
        RECT 10.650 4.260 11.050 6.880 ;
        RECT 10.450 4.850 11.050 6.880 ;
        RECT 10.450 1.040 11.050 1.490 ;
        RECT 10.650 1.040 11.050 1.920 ;
        RECT 9.670 0.840 10.070 1.490 ;
        RECT 9.720 2.400 11.230 2.700 ;
        RECT 10.830 2.320 11.230 2.720 ;
        RECT 9.720 0.840 10.020 6.670 ;
        RECT 9.670 4.850 10.070 6.670 ;
  END 
END NOR4X1

MACRO NOR3X1
  CLASS  CORE ;
  FOREIGN NOR3X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.920 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.940 1.400 1.340 1.800 ;
        RECT 0.770 1.500 1.340 1.800 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.450 2.110 1.850 2.980 ;
        RECT 2.700 2.630 3.100 3.030 ;
        RECT 1.450 2.680 3.100 2.980 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.410 1.450 6.420 1.850 ;
    END
  END C
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.740 -0.540 1.140 0.650 ;
        RECT 5.410 -0.540 7.010 0.650 ;
        RECT 0.000 -0.540 7.920 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.570 0.840 2.870 2.090 ;
        RECT 6.010 3.930 6.410 6.480 ;
        RECT 6.010 2.160 6.310 6.480 ;
        RECT 4.150 2.160 6.310 2.460 ;
        RECT 4.080 0.840 4.480 1.490 ;
        RECT 4.150 0.840 4.450 2.460 ;
        RECT 2.570 1.790 4.450 2.090 ;
        RECT 2.520 0.840 2.920 1.490 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.690 7.270 1.890 8.460 ;
        RECT 4.550 7.270 4.950 8.460 ;
        RECT 0.000 7.380 7.920 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 1.490 3.930 1.890 6.770 ;
        RECT 1.740 1.040 2.140 1.490 ;
        RECT 3.300 1.040 3.700 1.490 ;
        RECT 0.810 3.330 2.570 3.630 ;
        RECT 0.810 3.330 1.110 6.480 ;
        RECT 0.710 3.930 1.110 6.480 ;
        RECT 2.270 3.330 2.570 6.480 ;
        RECT 3.830 3.930 4.230 6.480 ;
        RECT 2.370 3.930 2.670 7.080 ;
        RECT 3.830 3.930 4.130 7.080 ;
        RECT 2.370 6.780 4.130 7.080 ;
        RECT 3.150 3.330 5.530 3.630 ;
        RECT 3.150 3.330 3.450 6.480 ;
        RECT 3.050 3.930 3.450 6.480 ;
        RECT 5.230 3.330 5.530 6.480 ;
        RECT 6.790 3.930 7.190 6.480 ;
        RECT 5.330 3.930 5.630 7.080 ;
        RECT 6.790 3.930 7.090 7.080 ;
        RECT 5.330 6.780 7.090 7.080 ;
  END 
END NOR3X1

MACRO NOR2X1
  CLASS  CORE ;
  FOREIGN NOR2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.300 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.750 2.770 1.150 3.830 ;
        RECT 0.750 3.430 1.180 3.830 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.110 2.110 2.630 2.510 ;
        RECT 2.230 2.110 2.630 2.840 ;
    END
  END B
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.670 -0.540 2.670 0.650 ;
        RECT 0.000 -0.540 3.300 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.510 1.250 1.810 3.770 ;
        RECT 2.230 4.070 2.630 6.670 ;
        RECT 2.230 3.470 2.530 6.670 ;
        RECT 1.510 3.470 2.530 3.770 ;
        RECT 1.450 2.770 1.850 3.170 ;
        RECT 1.450 1.250 1.850 1.900 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.670 7.270 2.690 8.460 ;
        RECT 0.000 7.380 3.300 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.670 4.510 1.070 6.770 ;
        RECT 0.670 1.150 1.070 1.900 ;
        RECT 1.450 4.070 1.850 6.670 ;
        RECT 2.230 1.150 2.630 1.780 ;
  END 
END NOR2X1

MACRO NAND4X1
  CLASS  CORE ;
  FOREIGN NAND4X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.430 3.040 3.830 3.830 ;
        RECT 3.430 3.040 4.140 3.440 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.770 4.090 3.170 4.860 ;
        RECT 2.770 4.460 3.360 4.860 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.110 3.040 2.510 3.830 ;
        RECT 2.110 3.040 2.580 3.440 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.790 4.090 1.190 4.860 ;
        RECT 0.790 4.460 1.680 4.860 ;
    END
  END D
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.540 5.280 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.880 5.260 2.280 7.080 ;
        RECT 1.880 5.260 4.840 5.660 ;
        RECT 4.440 2.240 4.840 5.660 ;
        RECT 4.220 0.840 4.620 2.640 ;
        RECT 4.090 4.090 4.840 4.490 ;
        RECT 3.440 5.260 3.840 7.080 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 7.380 5.280 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.500 5.260 1.500 6.880 ;
        RECT 0.500 1.040 1.500 2.640 ;
        RECT 1.880 0.840 2.280 2.640 ;
        RECT 2.660 6.210 3.060 6.880 ;
        RECT 2.660 0.840 3.060 2.640 ;
        RECT 3.440 0.840 3.840 2.640 ;
        RECT 4.220 6.210 4.620 6.880 ;
  END 
END NAND4X1

MACRO BUFX1
  CLASS  CORE ;
  FOREIGN BUFX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.960 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 2.820 1.800 3.240 ;
    END
  END A
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 -0.540 0.780 0.650 ;
        RECT 0.000 -0.540 3.960 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.110 4.270 2.410 6.670 ;
        RECT 2.110 4.270 3.120 4.570 ;
        RECT 2.820 2.440 3.120 4.570 ;
        RECT 2.460 0.840 2.860 2.740 ;
        RECT 2.060 4.870 2.460 6.670 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 7.270 3.300 8.460 ;
        RECT 0.000 7.380 3.960 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 1.280 4.870 1.680 6.770 ;
        RECT 1.280 1.040 2.080 2.440 ;
        RECT 0.500 1.740 0.900 2.440 ;
        RECT 0.500 3.650 2.400 3.950 ;
        RECT 2.000 3.560 2.400 3.960 ;
        RECT 0.500 1.740 0.800 6.670 ;
        RECT 0.500 4.870 0.900 6.670 ;
        RECT 2.840 4.870 3.240 6.770 ;
  END 
END BUFX1

MACRO NAND3X1
  CLASS  CORE ;
  FOREIGN NAND3X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.620 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 3.080 3.390 3.480 3.790 ;
        RECT 3.080 3.480 3.780 3.780 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.840 2.820 2.580 3.120 ;
        RECT 2.180 2.740 2.580 3.140 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.840 4.050 1.680 4.450 ;
    END
  END C
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.540 4.620 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.980 4.250 2.280 6.670 ;
        RECT 1.980 4.250 4.430 4.550 ;
        RECT 4.130 2.640 4.430 4.550 ;
        RECT 3.440 2.640 4.430 2.940 ;
        RECT 3.440 4.850 3.840 6.670 ;
        RECT 3.440 0.840 3.840 2.940 ;
        RECT 3.500 4.250 3.800 6.670 ;
        RECT 2.820 4.140 3.120 4.550 ;
        RECT 1.880 4.850 2.280 6.670 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.840 7.270 4.040 8.460 ;
        RECT 0.000 7.380 4.620 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 1.100 4.850 1.500 6.770 ;
        RECT 0.500 1.040 1.500 2.340 ;
        RECT 1.880 0.840 2.280 2.340 ;
        RECT 2.660 4.850 3.060 6.770 ;
        RECT 2.660 0.840 3.060 2.340 ;
  END 
END NAND3X1

MACRO NAND2X2
  CLASS  CORE ;
  FOREIGN NAND2X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.620 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.160 3.410 2.860 3.810 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.840 3.430 1.810 3.830 ;
    END
  END B
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.540 4.620 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.390 4.250 1.690 6.670 ;
        RECT 1.390 4.250 3.780 4.550 ;
        RECT 3.480 2.340 3.780 4.550 ;
        RECT 2.850 2.340 3.780 2.640 ;
        RECT 2.850 4.850 3.250 6.670 ;
        RECT 2.850 0.840 3.250 2.640 ;
        RECT 2.900 4.250 3.200 6.670 ;
        RECT 1.290 4.850 1.690 6.670 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.240 7.270 4.040 8.460 ;
        RECT 0.000 7.380 4.620 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.510 4.850 0.910 6.770 ;
        RECT 0.510 4.850 0.740 6.880 ;
        RECT 0.690 1.040 1.690 2.340 ;
        RECT 2.070 4.850 2.470 6.770 ;
        RECT 2.070 0.840 2.470 2.340 ;
        RECT 3.630 4.850 4.030 6.770 ;
  END 
END NAND2X2

MACRO NAND2X1
  CLASS  CORE ;
  FOREIGN NAND2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.300 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.790 3.430 1.190 4.490 ;
        RECT 0.790 3.430 1.250 3.830 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.160 3.740 2.560 4.440 ;
    END
  END B
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.560 -0.540 2.690 0.650 ;
        RECT 0.000 -0.540 3.300 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.730 1.250 1.130 1.900 ;
        RECT 1.560 2.820 2.460 3.120 ;
        RECT 1.510 4.850 1.910 6.670 ;
        RECT 1.560 2.200 1.860 6.670 ;
        RECT 0.830 2.200 1.860 2.500 ;
        RECT 0.830 1.250 1.130 2.500 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.580 7.270 2.690 8.460 ;
        RECT 0.000 7.380 3.300 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.730 4.850 1.130 6.770 ;
        RECT 1.510 1.250 1.910 1.900 ;
        RECT 2.290 4.850 2.690 6.770 ;
        RECT 2.290 1.150 2.690 1.900 ;
  END 
END NAND2X1

MACRO AND2X1
  CLASS  CORE ;
  FOREIGN AND2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.960 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.690 4.050 1.090 4.450 ;
        RECT 0.790 4.090 1.190 4.490 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.760 2.670 2.460 3.120 ;
        RECT 2.090 2.760 2.510 3.170 ;
    END
  END B
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.850 -0.540 3.250 0.650 ;
        RECT 0.000 -0.540 3.960 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.110 4.090 2.510 4.550 ;
        RECT 3.380 1.600 3.680 5.150 ;
        RECT 3.020 4.850 3.420 6.670 ;
        RECT 2.110 4.250 3.680 4.550 ;
        RECT 3.020 1.250 3.420 1.900 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.680 7.270 3.250 8.460 ;
        RECT 0.000 7.380 3.960 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.680 4.850 1.080 6.770 ;
        RECT 1.460 1.250 1.860 1.900 ;
        RECT 2.240 4.850 2.640 6.770 ;
        RECT 2.240 1.150 2.640 1.900 ;
        RECT 0.680 1.250 1.080 1.900 ;
        RECT 0.780 1.250 1.080 3.730 ;
        RECT 0.780 3.430 1.810 3.730 ;
        RECT 1.510 3.490 3.080 3.790 ;
        RECT 2.680 3.440 3.080 3.840 ;
        RECT 1.510 3.430 1.810 6.670 ;
        RECT 1.460 4.850 1.860 6.670 ;
  END 
END AND2X1

MACRO INVX8
  CLASS  CORE ;
  FOREIGN INVX8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.600 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.110 2.770 2.860 3.170 ;
    END
  END A
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 -0.540 0.900 0.650 ;
        RECT 5.620 -0.540 6.020 0.650 ;
        RECT 0.000 -0.540 6.600 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.550 4.180 1.950 6.670 ;
        RECT 4.670 4.180 5.070 6.670 ;
        RECT 1.550 4.180 5.070 4.580 ;
        RECT 2.280 1.940 4.240 2.340 ;
        RECT 3.840 0.840 4.240 2.340 ;
        RECT 3.430 1.940 3.830 4.580 ;
        RECT 3.110 4.180 3.510 6.670 ;
        RECT 2.280 0.840 2.680 2.340 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.770 7.270 5.970 8.460 ;
        RECT 0.000 7.380 6.600 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.770 4.180 1.170 6.770 ;
        RECT 1.500 1.040 1.900 2.340 ;
        RECT 2.330 5.020 2.730 6.770 ;
        RECT 3.060 1.040 3.460 1.240 ;
        RECT 3.890 5.020 4.290 6.770 ;
        RECT 4.620 1.040 5.020 2.340 ;
        RECT 5.450 4.180 5.850 6.770 ;
  END 
END INVX8

MACRO INVX4
  CLASS  CORE ;
  FOREIGN INVX4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.960 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.840 2.770 2.080 3.170 ;
    END
  END A
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.540 3.960 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.760 3.570 1.060 6.660 ;
        RECT 2.380 2.770 3.170 3.170 ;
        RECT 2.280 4.170 2.680 6.660 ;
        RECT 2.380 0.840 2.680 6.660 ;
        RECT 0.760 3.570 2.680 3.870 ;
        RECT 2.280 0.840 2.680 2.340 ;
        RECT 0.720 4.170 1.120 6.660 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.910 7.270 3.460 8.460 ;
        RECT 0.000 7.380 3.960 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 1.500 4.170 1.900 6.770 ;
        RECT 0.900 1.040 1.900 2.340 ;
        RECT 3.060 4.170 3.460 6.770 ;
        RECT 3.060 1.040 3.460 2.340 ;
  END 
END INVX4

MACRO INVX2
  CLASS  CORE ;
  FOREIGN INVX2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.300 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.780 3.430 1.510 3.830 ;
    END
  END A
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.540 3.300 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.820 4.250 1.120 6.670 ;
        RECT 2.280 4.850 2.680 6.670 ;
        RECT 2.280 0.840 2.680 2.340 ;
        RECT 2.280 0.840 2.580 6.670 ;
        RECT 0.820 4.250 2.580 4.550 ;
        RECT 2.160 3.480 2.580 3.780 ;
        RECT 0.720 4.850 1.120 6.670 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 7.270 2.500 8.460 ;
        RECT 0.000 7.380 3.300 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 1.500 4.850 1.900 6.770 ;
        RECT 0.900 1.040 1.900 2.340 ;
  END 
END INVX2

MACRO INVX1
  CLASS  CORE ;
  FOREIGN INVX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.640 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.790 3.430 1.190 4.280 ;
        RECT 0.790 3.880 1.310 4.280 ;
    END
  END A
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.720 -0.540 1.920 0.650 ;
        RECT 0.000 -0.540 2.640 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.510 1.250 1.910 1.900 ;
        RECT 1.510 4.850 1.910 6.670 ;
        RECT 1.610 1.250 1.910 6.670 ;
        RECT 1.500 2.820 1.910 3.120 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.720 7.270 1.920 8.460 ;
        RECT 0.000 7.380 2.640 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.730 4.850 1.130 6.770 ;
        RECT 0.730 1.150 1.130 1.900 ;
  END 
END INVX1

MACRO SDFFSRX1
  CLASS  CORE ;
  FOREIGN SDFFSRX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.640 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 32.470 1.360 32.975 2.010 ;
        RECT 32.730 2.770 33.540 3.170 ;
        RECT 32.690 4.650 33.090 6.470 ;
        RECT 32.730 2.310 33.030 6.470 ;
        RECT 32.675 1.360 32.975 2.610 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 34.250 1.360 34.650 2.010 ;
        RECT 34.350 3.480 34.800 3.780 ;
        RECT 34.250 4.650 34.650 6.470 ;
        RECT 34.350 1.360 34.650 6.470 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 6.120 3.430 6.920 3.830 ;
        RECT 6.520 3.430 6.920 3.835 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.140 4.750 4.940 5.150 ;
        RECT 4.540 4.750 4.940 5.280 ;
    END
  END SE
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.185 -0.540 3.085 0.650 ;
        RECT 0.000 -0.540 35.645 0.540 ;
        RECT 29.810 -0.540 31.210 0.650 ;
        RECT 7.120 -0.540 14.020 0.650 ;
    END
  END GRND
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 26.940 4.150 27.340 4.550 ;
        RECT 27.240 4.140 27.540 4.440 ;
    END
  END RN
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 5.620 4.840 6.020 5.280 ;
        RECT 8.165 4.205 8.565 4.605 ;
        RECT 6.120 4.210 8.565 4.510 ;
        RECT 5.610 4.840 6.420 5.140 ;
        RECT 6.120 4.210 6.420 5.140 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.730 3.430 1.280 3.830 ;
    END
  END CK
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.965 7.270 2.865 8.460 ;
        RECT 0.000 7.380 35.640 8.460 ;
        RECT 32.460 7.270 34.360 8.460 ;
        RECT 23.160 7.270 25.060 8.460 ;
        RECT 13.850 7.270 15.960 8.460 ;
        RECT 5.845 7.270 8.800 8.460 ;
    END
  END POWR
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 16.775 3.310 17.175 3.710 ;
        RECT 23.050 4.125 23.450 4.525 ;
        RECT 20.940 4.320 23.315 4.620 ;
        RECT 20.940 3.700 21.240 4.620 ;
        RECT 18.000 3.700 21.240 4.000 ;
        RECT 16.775 3.410 18.350 3.710 ;
        RECT 17.950 3.700 21.240 3.820 ;
    END
  END SN
  OBS 
      LAYER Metal1 ;
        RECT 1.380 5.620 1.780 6.770 ;
        RECT 1.680 1.150 2.080 1.795 ;
        RECT 0.500 1.395 0.900 1.795 ;
        RECT 0.470 1.425 0.770 2.790 ;
        RECT 0.470 2.490 2.070 2.790 ;
        RECT 1.770 2.490 2.070 4.920 ;
        RECT 0.650 4.600 2.165 4.900 ;
        RECT 1.765 4.520 2.165 4.920 ;
        RECT 0.650 4.600 0.950 6.020 ;
        RECT 0.600 5.620 1.000 6.020 ;
        RECT 2.610 1.395 3.260 1.795 ;
        RECT 2.610 3.650 3.110 4.050 ;
        RECT 2.610 1.395 2.910 5.920 ;
        RECT 2.160 5.620 2.910 5.920 ;
        RECT 2.160 5.620 2.560 6.020 ;
        RECT 4.540 6.185 4.940 6.880 ;
        RECT 4.935 1.040 5.340 1.795 ;
        RECT 5.320 6.185 6.720 6.585 ;
        RECT 8.400 6.185 8.800 6.770 ;
        RECT 3.760 1.395 4.160 1.795 ;
        RECT 3.760 1.395 4.025 2.400 ;
        RECT 9.370 4.885 9.770 5.285 ;
        RECT 7.130 4.985 9.770 5.285 ;
        RECT 3.470 2.100 3.770 6.575 ;
        RECT 7.130 4.985 7.430 5.880 ;
        RECT 3.470 5.580 7.430 5.880 ;
        RECT 3.470 5.580 4.070 6.575 ;
        RECT 3.725 1.400 3.770 6.575 ;
        RECT 3.760 6.185 4.160 6.585 ;
        RECT 7.750 5.585 9.960 5.885 ;
        RECT 9.660 5.585 9.960 6.585 ;
        RECT 7.750 5.585 8.050 6.550 ;
        RECT 7.500 6.185 7.900 6.585 ;
        RECT 9.660 6.185 10.060 6.585 ;
        RECT 10.170 1.150 10.570 2.045 ;
        RECT 4.940 2.705 7.520 3.005 ;
        RECT 7.220 2.705 7.520 3.865 ;
        RECT 4.070 3.650 4.470 4.050 ;
        RECT 7.220 3.565 9.875 3.865 ;
        RECT 4.940 2.705 5.240 4.050 ;
        RECT 4.070 3.750 5.240 4.050 ;
        RECT 9.575 3.565 9.875 4.485 ;
        RECT 11.105 4.085 11.505 4.485 ;
        RECT 9.575 4.185 11.505 4.485 ;
        RECT 11.440 6.185 11.840 6.880 ;
        RECT 4.340 2.095 8.120 2.395 ;
        RECT 7.820 2.095 8.120 3.255 ;
        RECT 4.340 2.095 4.640 3.145 ;
        RECT 4.240 2.745 4.640 3.145 ;
        RECT 7.820 2.955 10.740 3.255 ;
        RECT 10.440 2.955 10.740 3.605 ;
        RECT 10.440 3.305 12.610 3.605 ;
        RECT 12.210 3.300 12.610 3.700 ;
        RECT 10.270 4.885 10.670 5.285 ;
        RECT 12.220 4.885 12.620 5.285 ;
        RECT 10.255 4.985 12.620 5.285 ;
        RECT 6.905 1.375 7.305 1.775 ;
        RECT 6.905 1.475 9.210 1.775 ;
        RECT 13.010 1.635 13.410 2.035 ;
        RECT 12.530 1.735 13.410 2.035 ;
        RECT 8.510 1.475 9.210 2.045 ;
        RECT 8.910 1.475 9.210 2.645 ;
        RECT 12.530 1.735 12.830 2.645 ;
        RECT 8.910 2.345 12.830 2.645 ;
        RECT 11.930 1.035 14.010 1.335 ;
        RECT 11.930 1.035 12.230 2.035 ;
        RECT 11.830 1.635 12.230 2.035 ;
        RECT 13.430 2.580 14.010 2.980 ;
        RECT 13.710 1.035 14.010 2.980 ;
        RECT 13.130 2.680 13.430 5.885 ;
        RECT 10.540 5.585 13.430 5.885 ;
        RECT 12.595 5.585 13.040 6.390 ;
        RECT 10.540 5.585 10.840 6.585 ;
        RECT 10.440 6.185 10.840 6.585 ;
        RECT 12.700 6.185 13.100 6.585 ;
        RECT 13.770 3.505 14.170 3.905 ;
        RECT 13.770 3.505 14.070 6.205 ;
        RECT 13.730 5.805 14.130 6.205 ;
        RECT 15.560 5.930 15.960 6.770 ;
        RECT 15.270 4.335 15.670 4.920 ;
        RECT 15.270 4.620 17.055 4.920 ;
        RECT 16.655 4.620 17.055 5.025 ;
        RECT 14.365 0.960 16.970 1.260 ;
        RECT 14.365 0.960 14.665 1.960 ;
        RECT 16.670 0.960 16.970 1.960 ;
        RECT 14.310 1.560 14.710 1.960 ;
        RECT 16.670 1.560 17.070 1.960 ;
        RECT 15.190 1.560 15.890 1.960 ;
        RECT 15.190 1.560 15.490 2.800 ;
        RECT 14.475 2.500 15.490 2.800 ;
        RECT 14.370 4.885 14.775 5.285 ;
        RECT 17.660 5.130 18.060 5.630 ;
        RECT 14.475 5.330 18.060 5.630 ;
        RECT 14.475 2.500 14.775 6.330 ;
        RECT 14.475 5.930 15.180 6.330 ;
        RECT 17.850 1.040 18.250 1.960 ;
        RECT 18.995 5.615 19.395 6.015 ;
        RECT 19.000 5.615 19.395 6.880 ;
        RECT 15.075 3.260 15.475 3.760 ;
        RECT 15.075 3.460 16.370 3.760 ;
        RECT 16.070 3.460 16.370 4.320 ;
        RECT 16.070 4.020 17.665 4.320 ;
        RECT 17.365 4.020 17.665 4.715 ;
        RECT 20.190 4.315 20.590 4.715 ;
        RECT 17.365 4.415 20.590 4.715 ;
        RECT 20.515 1.040 20.910 1.715 ;
        RECT 20.510 1.315 20.910 1.715 ;
        RECT 15.995 2.265 19.595 2.560 ;
        RECT 17.575 2.260 19.595 2.560 ;
        RECT 15.870 2.360 17.875 2.565 ;
        RECT 19.295 2.260 19.595 2.925 ;
        RECT 15.870 2.360 16.270 2.760 ;
        RECT 19.295 2.625 22.150 2.925 ;
        RECT 21.850 2.625 22.150 3.920 ;
        RECT 22.150 3.620 22.550 4.020 ;
        RECT 22.810 5.520 23.210 5.920 ;
        RECT 21.055 6.295 21.455 6.695 ;
        RECT 22.905 5.520 23.205 6.695 ;
        RECT 21.055 6.395 23.205 6.695 ;
        RECT 23.075 1.040 23.470 2.030 ;
        RECT 23.070 1.630 23.470 2.030 ;
        RECT 24.070 5.520 24.470 6.770 ;
        RECT 18.850 1.365 20.210 1.665 ;
        RECT 21.410 1.630 21.810 2.030 ;
        RECT 18.850 1.315 19.250 1.715 ;
        RECT 19.910 1.365 20.210 2.315 ;
        RECT 21.410 1.680 22.750 2.030 ;
        RECT 19.910 2.015 21.715 2.315 ;
        RECT 22.450 1.680 22.750 3.035 ;
        RECT 22.450 2.735 23.150 3.035 ;
        RECT 22.850 2.735 23.150 3.825 ;
        RECT 22.850 3.525 24.050 3.825 ;
        RECT 23.750 3.525 24.050 5.220 ;
        RECT 25.150 4.720 25.550 5.220 ;
        RECT 22.210 4.920 25.570 5.220 ;
        RECT 18.360 5.015 20.555 5.315 ;
        RECT 20.255 5.015 20.555 6.015 ;
        RECT 22.210 4.920 22.510 5.950 ;
        RECT 20.255 5.650 22.510 5.950 ;
        RECT 20.255 5.615 20.655 6.015 ;
        RECT 16.820 5.930 17.220 6.330 ;
        RECT 18.360 5.015 18.660 6.330 ;
        RECT 16.820 6.030 18.660 6.330 ;
        RECT 24.070 1.085 26.485 1.385 ;
        RECT 26.185 1.085 26.485 2.085 ;
        RECT 24.070 1.085 24.370 2.085 ;
        RECT 23.970 1.685 24.370 2.085 ;
        RECT 26.185 1.435 26.730 2.085 ;
        RECT 27.110 1.040 27.510 2.085 ;
        RECT 28.305 3.665 28.705 4.065 ;
        RECT 28.305 3.665 28.605 4.650 ;
        RECT 27.920 4.350 28.605 4.650 ;
        RECT 27.920 4.350 28.220 6.520 ;
        RECT 25.885 6.430 28.145 6.730 ;
        RECT 27.745 4.950 28.145 6.770 ;
        RECT 25.835 6.530 26.235 6.930 ;
        RECT 28.525 4.950 28.925 6.880 ;
        RECT 27.890 1.600 29.095 1.900 ;
        RECT 28.695 1.585 29.095 1.985 ;
        RECT 27.890 1.435 28.290 2.085 ;
        RECT 24.965 3.025 29.700 3.325 ;
        RECT 29.310 3.085 29.710 3.485 ;
        RECT 26.350 3.025 26.750 3.505 ;
        RECT 24.965 3.025 25.365 3.590 ;
        RECT 25.150 1.685 25.550 2.085 ;
        RECT 25.180 1.685 25.480 2.690 ;
        RECT 23.510 2.390 30.410 2.690 ;
        RECT 23.510 2.390 23.910 3.090 ;
        RECT 30.110 2.390 30.410 3.730 ;
        RECT 30.030 3.430 31.190 3.730 ;
        RECT 30.790 3.400 31.190 3.800 ;
        RECT 24.360 2.390 24.660 4.220 ;
        RECT 24.360 3.920 26.320 4.220 ;
        RECT 30.030 3.430 30.330 6.395 ;
        RECT 26.020 3.920 26.320 5.820 ;
        RECT 25.330 5.520 26.320 5.820 ;
        RECT 25.330 5.520 25.730 5.920 ;
        RECT 29.930 5.695 30.330 6.395 ;
        RECT 30.910 5.245 31.310 6.880 ;
        RECT 30.910 6.240 31.315 6.880 ;
        RECT 31.710 1.040 32.090 2.010 ;
        RECT 31.690 1.150 32.090 2.010 ;
        RECT 30.510 1.345 31.035 1.745 ;
        RECT 30.735 1.345 31.035 2.640 ;
        RECT 30.735 2.340 32.255 2.640 ;
        RECT 31.870 2.410 32.270 2.810 ;
        RECT 31.890 3.880 32.290 4.280 ;
        RECT 31.955 2.340 32.255 4.545 ;
        RECT 31.735 4.245 32.035 6.395 ;
        RECT 31.690 5.245 32.090 6.395 ;
        RECT 33.470 4.650 33.870 6.770 ;
        RECT 33.470 1.040 33.870 2.010 ;
  END 
END SDFFSRX1

MACRO BUF_INVX8
  CLASS  CORE ;
  FOREIGN BUF_INVX8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.600 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.110 2.770 2.860 3.170 ;
    END
  END A
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 -0.540 0.900 0.650 ;
        RECT 5.620 -0.540 6.020 0.650 ;
        RECT 0.000 -0.540 6.600 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.550 4.180 1.950 6.670 ;
        RECT 4.670 4.180 5.070 6.670 ;
        RECT 1.550 4.180 5.070 4.580 ;
        RECT 2.280 1.940 4.240 2.340 ;
        RECT 3.840 0.840 4.240 2.340 ;
        RECT 3.430 1.940 3.830 4.580 ;
        RECT 3.110 4.180 3.510 6.670 ;
        RECT 2.280 0.840 2.680 2.340 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.770 7.270 5.970 8.460 ;
        RECT 0.000 7.380 6.600 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.770 4.180 1.170 6.770 ;
        RECT 1.500 1.040 1.900 2.340 ;
        RECT 2.330 5.020 2.730 6.770 ;
        RECT 3.060 1.040 3.460 1.240 ;
        RECT 3.890 5.020 4.290 6.770 ;
        RECT 4.620 1.040 5.020 2.340 ;
        RECT 5.450 4.180 5.850 6.770 ;
  END 
END BUF_INVX8

MACRO BUF_INVX4
  CLASS  CORE ;
  FOREIGN BUF_INVX4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.960 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.840 2.770 2.080 3.170 ;
    END
  END A
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.540 3.960 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.760 3.570 1.060 6.660 ;
        RECT 2.380 2.770 3.170 3.170 ;
        RECT 2.280 4.170 2.680 6.660 ;
        RECT 2.380 0.840 2.680 6.660 ;
        RECT 0.760 3.570 2.680 3.870 ;
        RECT 2.280 0.840 2.680 2.340 ;
        RECT 0.720 4.170 1.120 6.660 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.910 7.270 3.460 8.460 ;
        RECT 0.000 7.380 3.960 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 1.500 4.170 1.900 6.770 ;
        RECT 0.900 1.040 1.900 2.340 ;
        RECT 3.060 4.170 3.460 6.770 ;
        RECT 3.060 1.040 3.460 2.340 ;
  END 
END BUF_INVX4

MACRO BUF_ITL
  CLASS  CORE ;
  FOREIGN BUF_ITL 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.300 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.780 3.430 1.510 3.830 ;
    END
  END A
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.540 3.300 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.820 4.250 1.120 6.670 ;
        RECT 2.280 4.850 2.680 6.670 ;
        RECT 2.280 0.840 2.680 2.340 ;
        RECT 2.280 0.840 2.580 6.670 ;
        RECT 0.820 4.250 2.580 4.550 ;
        RECT 2.160 3.480 2.580 3.780 ;
        RECT 0.720 4.850 1.120 6.670 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 7.270 2.500 8.460 ;
        RECT 0.000 7.380 3.300 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 1.500 4.850 1.900 6.770 ;
        RECT 0.900 1.040 1.900 2.340 ;
  END 
END BUF_ITL

MACRO BUF_INVX1
  CLASS  CORE ;
  FOREIGN BUF_INVX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.640 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.790 3.430 1.190 4.280 ;
        RECT 0.790 3.880 1.310 4.280 ;
    END
  END A
  PIN GRND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.720 -0.540 1.920 0.650 ;
        RECT 0.000 -0.540 2.640 0.540 ;
    END
  END GRND
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.510 1.250 1.910 1.900 ;
        RECT 1.510 4.850 1.910 6.670 ;
        RECT 1.610 1.250 1.910 6.670 ;
        RECT 1.500 2.820 1.910 3.120 ;
    END
  END Y
  PIN POWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.720 7.270 1.920 8.460 ;
        RECT 0.000 7.380 2.640 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 0.730 4.850 1.130 6.770 ;
        RECT 0.730 1.150 1.130 1.900 ;
  END 
END BUF_INVX1


END LIBRARY
