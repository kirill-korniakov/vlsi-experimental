# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2008, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use.  This file contains valuable trade secrets and    *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *           NGLibraryCreator Development_version build 0810081030            *
# *                                                                            *
# ******************************************************************************
# 
# 

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.0025 ;

LAYER metal1
  TYPE ROUTING ;
  WIDTH 0.065 ;
  SPACING 0.065 ;
  PITCH 0.19 0.14 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.38 ;
  THICKNESS 0.13 ;
  CAPACITANCE CPERSQDIST 7.71613e-05 ;
  EDGECAPACITANCE 3.86e-05 ;
END metal1

LAYER via1
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.065 ;
END via1

LAYER metal2
  TYPE ROUTING ;
  WIDTH 0.07 ;
  SPACING 0.07 ;
  PITCH 0.19 0.14 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.25 ;
  THICKNESS 0.14 ;
  CAPACITANCE CPERSQDIST 4.08957e-05 ;
  EDGECAPACITANCE 2.04e-05 ;
END metal2

LAYER via2
  TYPE CUT ;
  SPACING 0.085 ;
  WIDTH 0.07 ;
END via2

LAYER metal3
  TYPE ROUTING ;
  WIDTH 0.07 ;
  SPACING 0.07 ;
  PITCH 0.19 0.14 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.25 ;
  THICKNESS 0.14 ;
  CAPACITANCE CPERSQDIST 2.7745e-05 ;
  EDGECAPACITANCE 1.39e-05 ;
END metal3

LAYER via3
  TYPE CUT ;
  SPACING 0.085 ;
  WIDTH 0.07 ;
END via3

LAYER metal4
  TYPE ROUTING ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  PITCH 0.28 0.28 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  CAPACITANCE CPERSQDIST 2.07429e-05 ;
  EDGECAPACITANCE 1.04e-05 ;
END metal4

LAYER via4
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
END via4

LAYER metal5
  TYPE ROUTING ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  PITCH 0.28 0.28 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  CAPACITANCE CPERSQDIST 1.3527e-05 ;
  EDGECAPACITANCE 6.76e-06 ;
END metal5

LAYER via5
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
END via5

LAYER metal6
  TYPE ROUTING ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  PITCH 0.28 0.28 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  CAPACITANCE CPERSQDIST 1.00359e-05 ;
  EDGECAPACITANCE 5.02e-06 ;
END metal6

LAYER via6
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
END via6

LAYER metal7
  TYPE ROUTING ;
  WIDTH 0.4 ;
  SPACING 0.4 ;
  PITCH 0.8 0.8 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.075 ;
  THICKNESS 0.8 ;
  CAPACITANCE CPERSQDIST 7.97709e-06 ;
  EDGECAPACITANCE 3.99e-06 ;
END metal7

LAYER via7
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
END via7

LAYER metal8
  TYPE ROUTING ;
  WIDTH 0.4 ;
  SPACING 0.4 ;
  PITCH 0.8 0.8 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.075 ;
  THICKNESS 0.8 ;
  CAPACITANCE CPERSQDIST 5.0391e-06 ;
  EDGECAPACITANCE 2.52e-06 ;
END metal8

LAYER via8
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
END via8

LAYER metal9
  TYPE ROUTING ;
  WIDTH 0.8 ;
  SPACING 0.8 ;
  PITCH 1.6 1.6 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.03 ;
  THICKNESS 2 ;
  CAPACITANCE CPERSQDIST 3.68273e-06 ;
  EDGECAPACITANCE 1.84e-06 ;
END metal9

LAYER via9
  TYPE CUT ;
  SPACING 0.88 ;
  WIDTH 0.8 ;
END via9

LAYER metal10
  TYPE ROUTING ;
  WIDTH 0.8 ;
  SPACING 0.8 ;
  PITCH 1.6 1.6 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.03 ;
  THICKNESS 2 ;
  CAPACITANCE CPERSQDIST 2.21236e-06 ;
  EDGECAPACITANCE 1.11e-06 ;
END metal10

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA via1_0 DEFAULT
  RESISTANCE 6 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal1 ;
    RECT -0.0675 -0.0675 0.0675 0.0675 ;
  LAYER metal2 ;
    RECT -0.0675 -0.0675 0.0675 0.0675 ;
END via1_0

VIA via1_1 DEFAULT
  RESISTANCE 6 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal1 ;
    RECT -0.0675 -0.0675 0.0675 0.0675 ;
  LAYER metal2 ;
    RECT -0.035 -0.0675 0.035 0.0675 ;
END via1_1

VIA via1_2 DEFAULT
  RESISTANCE 6 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal1 ;
    RECT -0.0675 -0.0675 0.0675 0.0675 ;
  LAYER metal2 ;
    RECT -0.0675 -0.035 0.0675 0.035 ;
END via1_2

VIA via1_3 DEFAULT
  RESISTANCE 6 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal1 ;
    RECT -0.0325 -0.0675 0.0325 0.0675 ;
  LAYER metal2 ;
    RECT -0.0675 -0.0675 0.0675 0.0675 ;
END via1_3

VIA via1_4 DEFAULT
  RESISTANCE 6 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal1 ;
    RECT -0.0325 -0.0675 0.0325 0.0675 ;
  LAYER metal2 ;
    RECT -0.035 -0.0675 0.035 0.0675 ;
END via1_4

VIA via1_5 DEFAULT
  RESISTANCE 6 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal1 ;
    RECT -0.0325 -0.0675 0.0325 0.0675 ;
  LAYER metal2 ;
    RECT -0.0675 -0.035 0.0675 0.035 ;
END via1_5

VIA via1_6 DEFAULT
  RESISTANCE 6 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal1 ;
    RECT -0.0675 -0.0325 0.0675 0.0325 ;
  LAYER metal2 ;
    RECT -0.0675 -0.0675 0.0675 0.0675 ;
END via1_6

VIA via1_7 DEFAULT
  RESISTANCE 6 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal1 ;
    RECT -0.0675 -0.0325 0.0675 0.0325 ;
  LAYER metal2 ;
    RECT -0.035 -0.0675 0.035 0.0675 ;
END via1_7

VIA via1_8 DEFAULT
  RESISTANCE 6 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal1 ;
    RECT -0.0675 -0.0325 0.0675 0.0325 ;
  LAYER metal2 ;
    RECT -0.0675 -0.035 0.0675 0.035 ;
END via1_8

VIA via2_0 DEFAULT
  RESISTANCE 5 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2_0

VIA via2_1 DEFAULT
  RESISTANCE 5 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via2_1

VIA via2_2 DEFAULT
  RESISTANCE 5 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via2_2

VIA via2_3 DEFAULT
  RESISTANCE 5 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER metal3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2_3

VIA via2_4 DEFAULT
  RESISTANCE 5 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via2_4

VIA via2_5 DEFAULT
  RESISTANCE 5 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via2_5

VIA via2_6 DEFAULT
  RESISTANCE 5 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2_6

VIA via2_7 DEFAULT
  RESISTANCE 5 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via2_7

VIA via2_8 DEFAULT
  RESISTANCE 5 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via2_8

VIA via3_0 DEFAULT
  RESISTANCE 5 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3_0

VIA via3_1 DEFAULT
  RESISTANCE 5 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3_1

VIA via3_2 DEFAULT
  RESISTANCE 5 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3_2

VIA via4_0 DEFAULT
  RESISTANCE 3 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via4_0

VIA via5_0 DEFAULT
  RESISTANCE 3 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via5_0

VIA via6_0 DEFAULT
  RESISTANCE 3 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END via6_0

VIA via7_0 DEFAULT
  RESISTANCE 1 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END via7_0

VIA via8_0 DEFAULT
  RESISTANCE 1 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END via8_0

VIA via9_0 DEFAULT
  RESISTANCE 0.5 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER metal9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER metal10 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END via9_0

VIARULE Via1Array-0 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0.035 0.035 ;
     WIDTH 0.135 TO 1.4 ;
  LAYER metal2 ;
    ENCLOSURE 0.035 0.035 ;
     WIDTH 0.135 TO 1.4 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
    SPACING 0.14 BY 0.14 ;
END Via1Array-0

VIARULE Via2Array-0 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0.035 0.035 ;
     WIDTH 0.14 TO 1.55 ;
  LAYER metal3 ;
    ENCLOSURE 0.035 0.035 ;
     WIDTH 0.14 TO 1.55 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END Via2Array-0

VIARULE Via3Array-0 GENERATE
  LAYER metal3 ;
    ENCLOSURE 0.035 0.035 ;
     WIDTH 0.14 TO 1.55 ;
  LAYER metal4 ;
    ENCLOSURE 0.035 0.035 ;
     WIDTH 0.14 TO 1.55 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END Via3Array-0

VIARULE Via4Array-0 GENERATE
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via4Array-0

VIARULE Via5Array-0 GENERATE
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via5Array-0

VIARULE Via6Array-0 GENERATE
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER metal7 ;
    ENCLOSURE 0.13 0.13 ;
     WIDTH 0.4 TO 3 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via6Array-0

VIARULE Via7Array-0 GENERATE
  LAYER metal7 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.4 TO 8.4 ;
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.4 TO 8.4 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END Via7Array-0

VIARULE Via8Array-0 GENERATE
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.4 TO 8.4 ;
  LAYER metal9 ;
    ENCLOSURE 0.2 0.2 ;
     WIDTH 0.8 TO 8.4 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END Via8Array-0

VIARULE Via9Array-0 GENERATE
  LAYER metal10 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.8 TO 16.8 ;
  LAYER metal9 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.8 TO 16.8 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
    SPACING 1.68 BY 1.68 ;
END Via9Array-0

VIARULE Via1Array-1 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
     WIDTH 0.135 TO 1.4 ;
  LAYER metal2 ;
    ENCLOSURE 0.0025 0.035 ;
     WIDTH 0.135 TO 1.4 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
    SPACING 0.14 BY 0.14 ;
END Via1Array-1

VIARULE Via2Array-1 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
     WIDTH 0.14 TO 1.55 ;
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
     WIDTH 0.14 TO 1.55 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END Via2Array-1

VIARULE Via3Array-1 GENERATE
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
     WIDTH 0.14 TO 1.55 ;
  LAYER metal4 ;
    ENCLOSURE 0.035 0.035 ;
     WIDTH 0.14 TO 1.55 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END Via3Array-1

VIARULE Via4Array-1 GENERATE
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via4Array-1

VIARULE Via5Array-1 GENERATE
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via5Array-1

VIARULE Via6Array-1 GENERATE
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER metal7 ;
    ENCLOSURE 0.13 0.13 ;
     WIDTH 0.4 TO 3 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via6Array-1

VIARULE Via7Array-1 GENERATE
  LAYER metal7 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.4 TO 8.4 ;
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.4 TO 8.4 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END Via7Array-1

VIARULE Via8Array-1 GENERATE
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.4 TO 8.4 ;
  LAYER metal9 ;
    ENCLOSURE 0.2 0.2 ;
     WIDTH 0.8 TO 8.4 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END Via8Array-1

VIARULE Via9Array-1 GENERATE
  LAYER metal10 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.8 TO 16.8 ;
  LAYER metal9 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.8 TO 16.8 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
    SPACING 1.68 BY 1.68 ;
END Via9Array-1

VIARULE Via1Array-2 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
     WIDTH 0.135 TO 1.4 ;
  LAYER metal2 ;
    ENCLOSURE 0.035 0.0025 ;
     WIDTH 0.135 TO 1.4 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
    SPACING 0.14 BY 0.14 ;
END Via1Array-2

VIARULE Via2Array-2 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
     WIDTH 0.14 TO 1.55 ;
  LAYER metal3 ;
    ENCLOSURE 0.035 0 ;
     WIDTH 0.14 TO 1.55 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END Via2Array-2

VIARULE Via3Array-2 GENERATE
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
     WIDTH 0.14 TO 1.55 ;
  LAYER metal4 ;
    ENCLOSURE 0.035 0.035 ;
     WIDTH 0.14 TO 1.55 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END Via3Array-2

VIARULE Via4Array-2 GENERATE
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via4Array-2

VIARULE Via5Array-2 GENERATE
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via5Array-2

VIARULE Via6Array-2 GENERATE
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER metal7 ;
    ENCLOSURE 0.13 0.13 ;
     WIDTH 0.4 TO 3 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via6Array-2

VIARULE Via7Array-2 GENERATE
  LAYER metal7 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.4 TO 8.4 ;
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.4 TO 8.4 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END Via7Array-2

VIARULE Via8Array-2 GENERATE
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.4 TO 8.4 ;
  LAYER metal9 ;
    ENCLOSURE 0.2 0.2 ;
     WIDTH 0.8 TO 8.4 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END Via8Array-2

VIARULE Via9Array-2 GENERATE
  LAYER metal10 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.8 TO 16.8 ;
  LAYER metal9 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.8 TO 16.8 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
    SPACING 1.68 BY 1.68 ;
END Via9Array-2

VIARULE Via1Array-3 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0.035 0 ;
     WIDTH 0.135 TO 1.4 ;
  LAYER metal2 ;
    ENCLOSURE 0.0025 0.035 ;
     WIDTH 0.135 TO 1.4 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
    SPACING 0.14 BY 0.14 ;
END Via1Array-3

VIARULE Via2Array-3 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0.035 0 ;
     WIDTH 0.14 TO 1.55 ;
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
     WIDTH 0.14 TO 1.55 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END Via2Array-3

VIARULE Via3Array-3 GENERATE
  LAYER metal3 ;
    ENCLOSURE 0.035 0 ;
     WIDTH 0.14 TO 1.55 ;
  LAYER metal4 ;
    ENCLOSURE 0.035 0.035 ;
     WIDTH 0.14 TO 1.55 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END Via3Array-3

VIARULE Via4Array-3 GENERATE
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via4Array-3

VIARULE Via5Array-3 GENERATE
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via5Array-3

VIARULE Via6Array-3 GENERATE
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.14 TO 3 ;
  LAYER metal7 ;
    ENCLOSURE 0.13 0.13 ;
     WIDTH 0.4 TO 3 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via6Array-3

VIARULE Via7Array-3 GENERATE
  LAYER metal7 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.4 TO 8.4 ;
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.4 TO 8.4 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END Via7Array-3

VIARULE Via8Array-3 GENERATE
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.4 TO 8.4 ;
  LAYER metal9 ;
    ENCLOSURE 0.2 0.2 ;
     WIDTH 0.8 TO 8.4 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END Via8Array-3

VIARULE Via9Array-3 GENERATE
  LAYER metal10 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.8 TO 16.8 ;
  LAYER metal9 ;
    ENCLOSURE 0 0 ;
     WIDTH 0.8 TO 16.8 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
    SPACING 1.68 BY 1.68 ;
END Via9Array-3

SPACING
  SAMENET metal1 metal1 0.065 ;
  SAMENET metal2 metal2 0.07 ;
  SAMENET metal3 metal3 0.07 ;
  SAMENET metal4 metal4 0.14 ;
  SAMENET metal5 metal5 0.14 ;
  SAMENET metal6 metal6 0.14 ;
  SAMENET metal7 metal7 0.4 ;
  SAMENET metal8 metal8 0.4 ;
  SAMENET metal9 metal9 0.8 ;
  SAMENET metal10 metal10 0.8 ;
  SAMENET via1 via1 0.075 ;
  SAMENET via2 via2 0.085 ;
  SAMENET via3 via3 0.085 ;
  SAMENET via4 via4 0.16 ;
  SAMENET via5 via5 0.16 ;
  SAMENET via6 via6 0.16 ;
  SAMENET via7 via7 0.44 ;
  SAMENET via8 via8 0.44 ;
  SAMENET via9 via9 0.88 ;
  SAMENET via1 via2 0.0 STACK ;
  SAMENET via2 via3 0.0 STACK ;
  SAMENET via3 via4 0.0 STACK ;
  SAMENET via4 via5 0.0 STACK ;
  SAMENET via5 via6 0.0 STACK ;
  SAMENET via6 via7 0.0 STACK ;
  SAMENET via7 via8 0.0 STACK ;
  SAMENET via8 via9 0.0 STACK ;
END SPACING

SITE NCSU_FreePDK_45nm
  SYMMETRY y ;
  CLASS core ;
  SIZE 0.19 BY 1.4 ;
END NCSU_FreePDK_45nm

MACRO AND2_X1
  CLASS core ;
  FOREIGN AND2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.0675 1.315 0.0675 1.0425 0.1325 1.0425 0.1325 1.315 0.4425 1.315 0.4425 1.0425 0.5075 1.0425 0.5075 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.4225 0.1275 0.4225 0.1275 0.5575 0.0625 0.5575  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.5075 0.085 0.5075 0.3975 0.4425 0.3975 0.4425 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4025 0.8425 0.5075 0.8425 0.5075 0.9775 0.4025 0.9775  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.2775 0.6975 0.2775 0.6975 1.1175 0.6325 1.1175  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.0675 0.2225 0.1325 0.2225 0.1325 0.2925 0.2275 0.2925 0.2275 0.315 0.3175 0.315 0.3175 0.7125 0.5025 0.7125 0.5025 0.6425 0.5675 0.6425 0.5675 0.7775 0.3175 0.7775 0.3175 1.1175 0.2525 1.1175 0.2525 0.38 0.1775 0.38 0.1775 0.3575 0.0675 0.3575  ;
  END
END AND2_X1

MACRO AND2_X2
  CLASS core ;
  FOREIGN AND2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.0525 1.315 0.0525 1.1475 0.1175 1.1475 0.1175 1.315 0.4475 1.315 0.4475 1.0075 0.5125 1.0075 0.5125 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.4225 0.1275 0.4225 0.1275 0.5575 0.0625 0.5575  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.5075 0.085 0.5075 0.3575 0.4425 0.3575 0.4425 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4025 0.8075 0.4425 0.8075 0.4425 0.7025 0.5075 0.7025 0.5075 0.8775 0.5425 0.8775 0.5425 0.9425 0.4025 0.9425  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.3275 0.6975 0.3275 0.6975 1.2275 0.6325 1.2275  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.0675 0.2225 0.1325 0.2225 0.1325 0.2925 0.1975 0.2925 0.1975 0.3025 0.3025 0.3025 0.3025 0.5025 0.5675 0.5025 0.5675 0.6375 0.5025 0.6375 0.5025 0.5675 0.3025 0.5675 0.3025 1.2225 0.2375 1.2225 0.2375 0.3675 0.1625 0.3675 0.1625 0.3575 0.0675 0.3575  ;
  END
END AND2_X2

MACRO AND2_X4
  CLASS core ;
  FOREIGN AND2_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.1275 0.11 1.1275 0.11 1.315 0.44 1.315 0.44 1.0675 0.505 1.0675 0.505 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.7025 0.1275 0.7025 0.1275 0.8375 0.0625 0.8375  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.505 0.085 0.505 0.3825 0.44 0.3825 0.44 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.36 0.6375 0.425 0.6375 0.425 0.7375 0.5425 0.7375 0.5425 0.8025 0.36 0.8025  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.8775 0.625 0.8775 0.625 0.2525 0.69 0.2525 0.69 1.0175 0.625 1.0175 0.625 0.9425 0.4075 0.9425  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.3925 0.11 0.3925 0.11 0.5075 0.56 0.5075 0.56 0.6525 0.495 0.6525 0.495 0.5725 0.295 0.5725 0.295 1.2025 0.23 1.2025 0.23 0.5725 0.06 0.5725 0.06 0.55 0.045 0.55  ;
  END
END AND2_X4

MACRO AND3_X1
  CLASS core ;
  FOREIGN AND3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.27 1.315 0.27 1.0675 0.335 1.0675 0.335 1.315 0.65 1.315 0.65 1.0675 0.715 1.0675 0.715 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.545 0.3975 0.61 0.3975 0.61 0.4575 0.7325 0.4575 0.7325 0.5325 0.545 0.5325  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.215 0.5275 0.28 0.5275 0.28 0.5975 0.3525 0.5975 0.3525 0.6625 0.215 0.6625  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.715 0.085 0.715 0.345 0.65 0.345 0.65 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.1775 0.42 0.1775 0.42 0.5325 0.355 0.5325 0.355 0.2425 0.2175 0.2425  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.5975 0.7375 0.84 0.7375 0.84 0.225 0.905 0.225 0.905 1.1425 0.84 1.1425 0.84 0.8025 0.5975 0.8025  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.085 0.2725 0.15 0.2725 0.15 0.9375 0.71 0.9375 0.71 0.8675 0.775 0.8675 0.775 1.0025 0.525 1.0025 0.525 1.1425 0.46 1.1425 0.46 1.0025 0.15 1.0025 0.15 1.1425 0.085 1.1425  ;
  END
END AND3_X1

MACRO AND3_X2
  CLASS core ;
  FOREIGN AND3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 1.1375 0.295 1.1375 0.295 1.315 0.63 1.315 0.63 0.9975 0.695 0.9975 0.695 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.3175 0.585 0.3175 0.585 0.485 0.52 0.485 0.52 0.3825 0.4075 0.3825  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.19 0.4575 0.3525 0.4575 0.3525 0.5225 0.255 0.5225 0.255 0.5925 0.19 0.5925  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.69 0.085 0.69 0.265 0.625 0.265 0.625 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.33 0.6675 0.395 0.6675 0.395 0.7375 0.5425 0.7375 0.5425 0.8025 0.33 0.8025  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.5975 0.5975 0.815 0.5975 0.815 0.235 0.88 0.235 0.88 1.2175 0.815 1.2175 0.815 0.6625 0.5975 0.6625  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.895 0.06 0.895 0.06 0.225 0.125 0.225 0.125 0.8725 0.46 0.8725 0.46 0.8675 0.685 0.8675 0.685 0.7975 0.75 0.7975 0.75 0.9325 0.485 0.9325 0.485 1.2125 0.42 1.2125 0.42 0.9375 0.11 0.9375 0.11 1.2125 0.045 1.2125  ;
  END
END AND3_X2

MACRO AND3_X4
  CLASS core ;
  FOREIGN AND3_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2375 1.315 0.2375 1.1325 0.3025 1.1325 0.3025 1.315 0.6375 1.315 0.6375 0.9925 0.7025 0.9925 0.7025 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.5625 0.5375 0.5625 0.5375 0.6975 0.4425 0.6975  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1825 0.5275 0.2475 0.5275 0.2475 0.5975 0.3525 0.5975 0.3525 0.6625 0.1825 0.6625  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.7025 0.085 0.7025 0.4075 0.6375 0.4075 0.6375 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.1775 0.3875 0.1775 0.3875 0.4875 0.3225 0.4875 0.3225 0.2425 0.2175 0.2425  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.8225 0.2775 0.8875 0.2775 0.8875 0.9425 0.8225 0.9425  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.0525 0.2275 0.1175 0.2275 0.1175 1.0025 0.4275 1.0025 0.4275 0.8625 0.6925 0.8625 0.6925 0.5425 0.7575 0.5425 0.7575 0.9275 0.4925 0.9275 0.4925 1.2075 0.4275 1.2075 0.4275 1.0675 0.1175 1.0675 0.1175 1.2075 0.0525 1.2075  ;
  END
END AND3_X4

MACRO AND4_X1
  CLASS core ;
  FOREIGN AND4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.1375 0.11 1.1375 0.11 1.315 0.42 1.315 0.42 1.1375 0.485 1.1375 0.485 1.315 0.8 1.315 0.8 1.1375 0.865 1.1375 0.865 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.5975 0.505 0.5975 0.505 0.5275 0.57 0.5275 0.57 0.6625 0.4075 0.6625  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.8075 0.24 0.8075 0.24 0.8775 0.3525 0.8775 0.3525 0.9425 0.175 0.9425  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.865 0.085 0.865 0.345 0.8 0.345 0.8 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.1775 0.405 0.1775 0.405 0.5325 0.34 0.5325 0.34 0.2425 0.2175 0.2425  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.695 0.3975 0.76 0.3975 0.76 0.4575 0.9225 0.4575 0.9225 0.5325 0.695 0.5325  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.7875 0.7375 0.99 0.7375 0.99 0.225 1.055 0.225 1.055 1.2125 0.99 1.2125 0.99 0.8025 0.7875 0.8025  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.2725 0.11 0.2725 0.11 1.0075 0.86 1.0075 0.86 0.9375 0.925 0.9375 0.925 1.0725 0.675 1.0725 0.675 1.2125 0.61 1.2125 0.61 1.0725 0.295 1.0725 0.295 1.2125 0.23 1.2125 0.23 1.0725 0.045 1.0725  ;
  END
END AND4_X1

MACRO AND4_X2
  CLASS core ;
  FOREIGN AND4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.1375 0.11 1.1375 0.11 1.315 0.42 1.315 0.42 1.1375 0.485 1.1375 0.485 1.315 0.82 1.315 0.82 0.9975 0.885 0.9975 0.885 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.5975 0.52 0.5975 0.52 0.5275 0.585 0.5275 0.585 0.6625 0.4075 0.6625  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.19 0.8075 0.255 0.8075 0.255 0.8775 0.3525 0.8775 0.3525 0.9425 0.19 0.9425  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.88 0.085 0.88 0.2525 0.815 0.2525 0.815 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.1775 0.405 0.1775 0.405 0.5175 0.34 0.5175 0.34 0.2425 0.2175 0.2425  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.71 0.3175 0.9225 0.3175 0.9225 0.3825 0.775 0.3825 0.775 0.5175 0.71 0.5175  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.7875 0.5975 1.005 0.5975 1.005 0.2225 1.07 0.2225 1.07 1.2175 1.005 1.2175 1.005 0.6625 0.7875 0.6625  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.06 0.2575 0.125 0.2575 0.125 1.0075 0.61 1.0075 0.61 0.8675 0.875 0.8675 0.875 0.7975 0.94 0.7975 0.94 0.9325 0.675 0.9325 0.675 1.2125 0.61 1.2125 0.61 1.0725 0.295 1.0725 0.295 1.2125 0.23 1.2125 0.23 1.0725 0.06 1.0725  ;
  END
END AND4_X2

MACRO AND4_X4
  CLASS core ;
  FOREIGN AND4_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.1725 0.11 1.1725 0.11 1.315 0.42 1.315 0.42 1.1725 0.485 1.1725 0.485 1.315 0.82 1.315 0.82 1.0325 0.885 1.0325 0.885 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.7025 0.53 0.7025 0.53 0.8375 0.4425 0.8375  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.19 0.8425 0.3175 0.8425 0.3175 0.9775 0.19 0.9775  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.88 0.085 0.88 0.4075 0.815 0.4075 0.815 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.4225 0.405 0.4225 0.405 0.5575 0.2525 0.5575  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.4225 0.735 0.4225 0.735 0.5575 0.6325 0.5575  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.005 0.2775 1.07 0.2775 1.07 0.5625 1.0775 0.5625 1.0775 0.6975 1.07 0.6975 1.07 0.9825 1.005 0.9825  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.06 0.2725 0.125 0.2725 0.125 1.0425 0.61 1.0425 0.61 0.9025 0.875 0.9025 0.875 0.5825 0.94 0.5825 0.94 0.9675 0.675 0.9675 0.675 1.2475 0.61 1.2475 0.61 1.1075 0.295 1.1075 0.295 1.2475 0.23 1.2475 0.23 1.1075 0.06 1.1075  ;
  END
END AND4_X4

MACRO ANTENNA_X1
  CLASS core ;
  FOREIGN ANTENNA_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.19 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.15 0.1275 0.15 0.1275 1.25 0.0625 1.25  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.19 1.315 0.19 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.19 -0.085 0.19 0.085 0 0.085  ;
    END
  END VSS
END ANTENNA_X1

MACRO AOI211_X1
  CLASS core ;
  FOREIGN AOI211_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.8225 0.5625 0.8875 0.5625 0.8875 0.6975 0.8225 0.6975  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.8 1.315 0.8 1.3075 0.8 1.0825 0.8 0.89 0.865 0.89 0.865 1.0825 0.865 1.3075 0.865 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.71 0.085 0.71 0.235 0.575 0.235 0.575 0.085 0.11 0.085 0.11 0.23 0.045 0.23 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.4575 0.5425 0.4575 0.5425 0.5225 0.5325 0.5225 0.5325 0.6 0.4675 0.6 0.4675 0.5225 0.4075 0.5225  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.23 0.2825 0.3175 0.2825 0.3175 0.3025 0.42 0.3025 0.42 0.15 0.485 0.15 0.485 0.3025 0.8 0.3025 0.8 0.15 0.865 0.15 0.865 0.3675 0.8 0.3675 0.485 0.3675 0.3175 0.3675 0.3175 0.4175 0.295 0.4175 0.295 1.12 0.23 1.12 0.23 0.4175  ;
    END
  END ZN
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.4225 0.1275 0.4225 0.1275 0.5575 0.0625 0.5575  ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.36 0.69 0.425 0.69 0.425 0.7375 0.5425 0.7375 0.5425 0.8025 0.425 0.8025 0.425 0.825 0.36 0.825 0.36 0.8025 0.36 0.7375  ;
    END
  END C1
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.89 0.11 0.89 0.11 1.185 0.42 1.185 0.42 0.89 0.485 0.89 0.485 1.25 0.045 1.25  ;
  END
END AOI211_X1

MACRO AOI211_X2
  CLASS core ;
  FOREIGN AOI211_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.7325 0.4225 0.8875 0.4225 0.8875 0.5575 0.7325 0.5575  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.8225 1.315 0.8225 0.68 0.8875 0.68 0.8875 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.7125 0.085 0.7125 0.2275 0.6475 0.2275 0.6475 0.085 0.1325 0.085 0.1325 0.38 0.0675 0.38 0.0675 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.5925 0.535 0.6575 0.535 0.6575 0.7025 0.6975 0.7025 0.6975 0.8375 0.5925 0.8375  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.2825 0.4425 0.2825 0.4425 0.15 0.5075 0.15 0.5075 0.2925 0.8375 0.2925 0.8375 0.1975 0.9025 0.1975 0.9025 0.3575 0.5075 0.3575 0.5075 0.425 0.4425 0.425 0.4425 0.3475 0.3175 0.3475 0.3175 1.075 0.2525 1.075  ;
    END
  END ZN
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.535 0.1275 0.535 0.1275 0.6975 0.0625 0.6975  ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3825 0.535 0.4475 0.535 0.4475 0.5625 0.5075 0.5625 0.5075 0.6975 0.4425 0.6975 0.4425 0.67 0.3825 0.67  ;
    END
  END C1
  OBS
      LAYER metal1 ;
        POLYGON 0.0675 0.79 0.1325 0.79 0.1325 1.14 0.4425 1.14 0.4425 0.79 0.5075 0.79 0.5075 1.14 0.5075 1.205 0.4425 1.205 0.1325 1.205 0.0675 1.205 0.0675 1.14  ;
  END
END AOI211_X2

MACRO AOI211_X4
  CLASS core ;
  FOREIGN AOI211_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.71 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.2025 0.4225 1.2675 0.4225 1.2675 0.6275 1.2025 0.6275  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 1.18 1.315 1.18 1.035 1.245 1.035 1.245 1.315 1.71 1.315 1.71 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.71 -0.085 1.71 0.085 1.245 0.085 1.245 0.3575 1.18 0.3575 1.18 0.085 0.865 0.085 0.865 0.38 0.8 0.38 0.8 0.085 0.11 0.085 0.11 0.38 0.045 0.38 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.915 0.6025 0.98 0.6025 0.98 0.6925 1.455 0.6925 1.455 0.6025 1.52 0.6025 1.52 0.7575 1.0775 0.7575 1.0775 0.8375 1.0125 0.8375 1.0125 0.7575 0.915 0.7575  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.775 0.785 0.775 0.785 0.51 0.425 0.51 0.425 0.15 0.49 0.15 0.49 0.2825 0.5075 0.2825 0.5075 0.445 0.99 0.445 0.99 0.2275 1.055 0.2275 1.055 0.51 0.85 0.51 0.85 0.84 0.675 0.84 0.675 1.05 0.61 1.05 0.61 0.84 0.3 0.84 0.3 1.05 0.235 1.05  ;
    END
  END ZN
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.5625 0.215 0.5625 0.215 0.6325 0.655 0.6325 0.655 0.575 0.72 0.575 0.72 0.71 0.655 0.71 0.655 0.6975 0.0625 0.6975  ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.2825 0.345 0.2825 0.345 0.55 0.28 0.55 0.28 0.4175 0.2525 0.4175  ;
    END
  END C1
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.905 0.11 0.905 0.11 1.115 0.42 1.115 0.42 0.905 0.485 0.905 0.485 1.115 0.8 1.115 0.8 1.015 0.805 1.015 0.805 0.905 1.625 0.905 1.625 1.18 1.56 1.18 1.56 0.97 0.87 0.97 0.87 1.04 0.865 1.04 0.865 1.18 0.045 1.18  ;
  END
END AOI211_X4

MACRO AOI21_X1
  CLASS core ;
  FOREIGN AOI21_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.7275 0.57 0.7275 0.57 0.8625 0.505 0.8625 0.505 0.8025 0.4075 0.8025  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.61 1.315 0.61 0.975 0.675 0.975 0.675 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.1775 0.36 0.1775 0.36 0.5325 0.295 0.5325 0.295 0.2425 0.2175 0.2425  ;
    END
  END B1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.675 0.085 0.675 0.3925 0.61 0.3925 0.61 0.085 0.11 0.085 0.11 0.3525 0.045 0.3525 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.4225 0.1275 0.4225 0.1275 0.5575 0.0625 0.5575  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.605 0.2675 0.605 0.2675 0.5975 0.425 0.5975 0.425 0.2725 0.49 0.2725 0.49 0.5975 0.5425 0.5975 0.5425 0.6625 0.3 0.6625 0.3 0.9875 0.235 0.9875  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.975 0.11 0.975 0.11 1.0525 0.42 1.0525 0.42 0.975 0.485 0.975 0.485 1.1175 0.045 1.1175  ;
  END
END AOI21_X1

MACRO AOI21_X2
  CLASS core ;
  FOREIGN AOI21_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.5975 0.6975 0.5975 0.6975 0.8375 0.6325 0.8375  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.6475 1.315 0.6475 0.9025 0.7125 0.9025 0.7125 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.4225 0.3625 0.4225 0.3625 0.5575 0.2525 0.5575  ;
    END
  END B1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.7125 0.085 0.7125 0.2475 0.6475 0.2475 0.6475 0.085 0.1325 0.085 0.1325 0.3875 0.0675 0.3875 0.0675 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.5625 0.1275 0.5625 0.1275 0.6975 0.0625 0.6975  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2725 0.6425 0.3025 0.6425 0.3025 0.6325 0.4425 0.6325 0.4425 0.1575 0.5075 0.1575 0.5075 0.6975 0.3375 0.6975 0.3375 0.9975 0.2725 0.9975  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.0825 0.8525 0.1475 0.8525 0.1475 1.0625 0.4575 1.0625 0.4575 0.8525 0.5225 0.8525 0.5225 1.1275 0.0825 1.1275  ;
  END
END AOI21_X2

MACRO AOI21_X4
  CLASS core ;
  FOREIGN AOI21_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.0125 0.5625 1.0775 0.5625 1.0775 0.8375 1.0125 0.8375  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.98 1.315 0.98 1.0325 1.115 1.0325 1.115 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.18 0.585 0.8275 0.585 0.8275 0.65 0.7325 0.65 0.7325 0.6625 0.5975 0.6625 0.5975 0.65 0.18 0.65  ;
    END
  END B1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 1.115 0.085 1.115 0.2975 0.98 0.2975 0.98 0.085 0.545 0.085 0.545 0.39 0.41 0.39 0.41 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3375 0.715 0.5525 0.715 0.5525 0.8025 0.3375 0.8025  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.05 0.455 0.07 0.455 0.07 0.195 0.135 0.195 0.135 0.455 0.825 0.455 0.825 0.195 0.89 0.195 0.89 0.52 0.115 0.52 0.115 0.8775 0.635 0.8775 0.635 0.8175 0.7 0.8175 0.7 1.0925 0.635 1.0925 0.635 0.9425 0.32 0.9425 0.32 1.12 0.255 1.12 0.255 0.9425 0.05 0.9425  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.51 1.185 0.825 1.185 0.825 0.9025 1.27 0.9025 1.27 1.1775 1.205 1.1775 1.205 0.9675 0.89 0.9675 0.89 1.25 0.07 1.25 0.07 1.115 0.135 1.115 0.135 1.185 0.445 1.185 0.445 1.075 0.41 1.075 0.41 1.01 0.545 1.01 0.545 1.075 0.51 1.075  ;
  END
END AOI21_X4

MACRO AOI221_X1
  CLASS core ;
  FOREIGN AOI221_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.5975 0.485 0.5975 0.485 0.526 0.55 0.526 0.55 0.6625 0.4075 0.6625  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 0.8675 0.295 0.8675 0.295 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.4225 0.34 0.4225 0.34 0.5575 0.2525 0.5575  ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.42 0.1775 0.485 0.1775 0.485 0.3775 0.99 0.3775 0.99 0.1925 1.055 0.1925 1.055 0.2825 1.0775 0.2825 1.0775 0.4425 0.87 0.4425 0.87 1.0975 0.805 1.0975 0.805 0.4425 0.42 0.4425  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.935 0.5625 1.0775 0.5625 1.0775 0.6975 0.935 0.6975  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.675 0.085 0.675 0.3125 0.61 0.3125 0.61 0.085 0.11 0.085 0.11 0.2725 0.045 0.2725 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.4225 0.1275 0.4225 0.1275 0.5575 0.0625 0.5575  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.5625 0.74 0.5625 0.74 0.6975 0.6325 0.6975  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.7375 0.485 0.7375 0.485 1.0975 0.42 1.0975 0.42 0.8025 0.11 0.8025 0.11 1.0975 0.045 1.0975  ;
        POLYGON 0.615 0.8675 0.68 0.8675 0.68 1.1625 0.99 1.1625 0.99 0.8675 1.055 0.8675 1.055 1.2275 0.615 1.2275  ;
  END
END AOI221_X1

MACRO AOI221_X2
  CLASS core ;
  FOREIGN AOI221_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.4575 0.53 0.4575 0.63 0.4575 0.63 0.5225 0.53 0.5225 0.4075 0.5225  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 1.0075 0.295 1.0075 0.295 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.5625 0.34 0.5625 0.34 0.6975 0.2525 0.6975  ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.385 0.325 0.42 0.325 0.42 0.15 0.485 0.15 0.485 0.325 0.8875 0.325 0.8875 0.39 0.8875 0.4 1.02 0.4 1.02 0.15 1.085 0.15 1.085 0.465 0.8875 0.465 0.8875 0.975 0.8225 0.975 0.8225 0.39 0.485 0.39 0.42 0.39 0.385 0.39  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.0125 0.575 1.0775 0.575 1.0775 0.8375 1.0125 0.8375  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.71 0.085 0.71 0.24 0.645 0.24 0.645 0.085 0.11 0.085 0.11 0.38 0.045 0.38 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.5625 0.1275 0.5625 0.1275 0.6975 0.0625 0.6975  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.5975 0.5975 0.6925 0.5975 0.6925 0.575 0.7575 0.575 0.7575 0.71 0.6925 0.71 0.6925 0.6625 0.5975 0.6625  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.8775 0.485 0.8775 0.485 1.1525 0.42 1.1525 0.42 0.9425 0.11 0.9425 0.11 1.1525 0.045 1.1525  ;
        POLYGON 0.6325 0.9025 0.6975 0.9025 0.6975 1.1125 1.0075 1.1125 1.0075 0.9025 1.0725 0.9025 1.0725 1.1775 0.6325 1.1775  ;
  END
END AOI221_X2

MACRO AOI221_X4
  CLASS core ;
  FOREIGN AOI221_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.28 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.2025 0.5625 1.2675 0.5625 1.2675 0.6975 1.2025 0.6975  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 1.52 1.315 1.52 1.0475 1.585 1.0475 1.585 1.315 1.9 1.315 1.9 1.0475 1.965 1.0475 1.965 1.315 2.28 1.315 2.28 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.795 0.415 1.86 0.415 1.86 0.4575 2.2175 0.4575 2.2175 0.5575 2.1525 0.5575 2.1525 0.5225 1.86 0.5225 1.86 0.55 1.795 0.55  ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.045 0.7775 0.2525 0.7775 0.2525 0.15 0.34 0.15 0.34 0.41 1.03 0.41 1.03 0.15 1.095 0.15 1.095 0.41 1.645 0.41 1.645 0.15 1.71 0.15 1.71 0.475 0.3175 0.475 0.3175 0.7775 0.485 0.7775 0.485 0.9675 0.8 0.9675 0.8 0.8325 0.865 0.8325 0.865 1.1075 0.8 1.1075 0.8 1.0325 0.485 1.0325 0.485 1.0525 0.42 1.0525 0.42 0.8425 0.11 0.8425 0.11 1.0525 0.045 1.0525  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3825 0.54 0.85 0.54 0.85 0.5625 0.8875 0.5625 0.8875 0.6975 0.8225 0.6975 0.8225 0.675 0.785 0.675 0.785 0.605 0.3825 0.605  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.28 -0.085 2.28 0.085 2.09 0.085 2.09 0.38 2.025 0.38 2.025 0.085 1.365 0.085 1.365 0.345 1.23 0.345 1.23 0.085 0.75 0.085 0.75 0.345 0.615 0.345 0.615 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.415 0.5625 1.6475 0.5625 1.6475 0.615 2.01 0.615 2.01 0.75 1.945 0.75 1.945 0.6975 1.415 0.6975  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.535 0.67 0.5975 0.67 0.67 0.67 0.67 0.7375 0.7325 0.7375 0.7325 0.8025 0.5975 0.8025 0.5975 0.7375 0.5975 0.735 0.535 0.735  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.235 0.9075 0.3 0.9075 0.3 1.1175 0.61 1.1175 0.61 1.1025 0.675 1.1025 0.675 1.1725 1.14 1.1725 1.14 0.9625 1.205 0.9625 1.205 1.2375 0.61 1.2375 0.61 1.1825 0.235 1.1825  ;
        POLYGON 0.955 0.8325 1.33 0.8325 1.33 0.76 1.395 0.76 1.395 0.8725 1.715 0.8725 1.715 0.7625 1.78 0.7625 1.78 0.8325 2.09 0.8325 2.09 0.74 2.155 0.74 2.155 1.015 2.09 1.015 2.09 0.8975 1.775 0.8975 1.775 1.0375 1.71 1.0375 1.71 0.9375 1.4 0.9375 1.4 1.035 1.335 1.035 1.335 0.8975 1.02 0.8975 1.02 1.1075 0.955 1.1075  ;
  END
END AOI221_X4

MACRO AOI222_X1
  CLASS core ;
  FOREIGN AOI222_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.5225 1.315 0.5225 1.055 0.5875 1.055 0.5875 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.7825 0.52 0.8225 0.52 0.825 0.52 0.8875 0.52 0.9175 0.52 0.9175 0.585 0.8875 0.585 0.8875 0.6975 0.8225 0.6975 0.8225 0.585 0.7825 0.585  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.0125 0.45 1.1275 0.45 1.1275 0.5625 1.1275 0.585 1.0775 0.585 1.0775 0.6975 1.0125 0.6975 1.0125 0.5625  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.3925 0.5625 1.4575 0.5625 1.4575 0.6975 1.3925 0.6975  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.1325 0.905 1.2025 0.905 1.2025 0.385 0.9875 0.385 0.9875 0.215 0.7425 0.215 0.7425 0.325 0.5975 0.325 0.5975 0.1775 0.6875 0.1775 0.6875 0.15 1.0525 0.15 1.0525 0.32 1.2675 0.32 1.2675 1.11 1.1325 1.11  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.5375 0.52 0.6325 0.52 0.635 0.52 0.6975 0.52 0.6975 0.6975 0.6325 0.6975 0.6325 0.585 0.5375 0.585  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 1.4275 0.085 1.4275 0.385 1.3625 0.385 1.3625 0.085 0.3625 0.085 0.3625 0.325 0.2275 0.325 0.2275 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.045 0.52 0.0625 0.52 0.0775 0.52 0.1425 0.52 0.18 0.52 0.18 0.585 0.1425 0.585 0.1275 0.585 0.1275 0.6975 0.0625 0.6975 0.0625 0.585 0.045 0.585  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.52 0.3175 0.52 0.4725 0.52 0.4725 0.585 0.3175 0.585 0.3175 0.6975 0.2525 0.6975  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.2975 0.91 0.8075 0.91 0.8075 1.115 0.6525 1.115 0.6525 0.975 0.4575 0.975 0.4575 1.115 0.2975 1.115  ;
        POLYGON 0.0775 0.28 0.1425 0.28 0.1425 0.39 0.8325 0.39 0.8325 0.28 0.8975 0.28 0.8975 0.415 0.8925 0.415 0.8925 0.455 0.0775 0.455  ;
        POLYGON 0.0625 0.78 1.0475 0.78 1.0475 1.175 1.3575 1.175 1.3575 0.915 1.4225 0.915 1.4225 1.24 0.9825 1.24 0.9825 0.845 0.1275 0.845 0.1275 0.91 0.1875 0.91 0.1875 1.185 0.0625 1.185  ;
  END
END AOI222_X1

MACRO AOI222_X2
  CLASS core ;
  FOREIGN AOI222_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.71 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.5175 1.315 0.5175 1.0675 0.5825 1.0675 0.5825 1.315 1.71 1.315 1.71 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6975 0.67 0.8225 0.67 0.8225 0.5625 0.8875 0.5625 0.8875 0.735 0.8525 0.735 0.8225 0.735 0.6975 0.735  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.0125 0.4225 1.165 0.4225 1.165 0.495 1.0775 0.495 1.0775 0.5575 1.0125 0.5575 1.0125 0.495 1.0125 0.49  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.36 0.5625 1.4575 0.5625 1.4575 0.6975 1.36 0.6975  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.2025 0.7025 1.23 0.7025 1.23 0.355 1.01 0.355 1.01 0.215 0.6125 0.215 0.6125 0.15 1.145 0.15 1.145 0.29 1.295 0.29 1.295 0.7025 1.295 0.8375 1.295 1.035 1.23 1.035 1.23 0.8375 1.2025 0.8375  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.5625 0.41 0.6975 0.41 0.6975 0.475 0.6975 0.5575 0.6325 0.5575 0.6325 0.475 0.5625 0.475  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.71 -0.085 1.71 0.085 1.53 0.085 1.53 0.36 1.465 0.36 1.465 0.085 0.3625 0.085 0.3625 0.165 0.2275 0.165 0.2275 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.5625 0.3175 0.5625 0.3175 0.6975 0.2525 0.6975  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.5625 0.5075 0.5625 0.5075 0.6975 0.4425 0.6975  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.3325 0.9375 0.7725 0.9375 0.7725 1.2125 0.7075 1.2125 0.7075 1.0025 0.3975 1.0025 0.3975 1.2125 0.3325 1.2125  ;
        POLYGON 0.0425 0.28 0.9325 0.28 0.9325 0.345 0.0425 0.345  ;
        POLYGON 0.125 0.8075 0.19 0.8075 0.9175 0.8075 0.9825 0.8075 0.9825 0.8725 0.9825 1.0425 0.9825 1.1 1.415 1.1 1.415 0.89 1.48 0.89 1.48 1.165 0.9175 1.165 0.9175 1.1 0.9175 1.0425 0.9175 0.8725 0.19 0.8725 0.19 0.97 0.19 1.14 0.125 1.14 0.125 0.97 0.125 0.8725  ;
  END
END AOI222_X2

MACRO AOI222_X4
  CLASS core ;
  FOREIGN AOI222_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.66 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 1.0325 0.295 1.0325 0.295 1.315 0.61 1.315 0.61 1.0325 0.675 1.0325 0.675 1.315 2.66 1.315 2.66 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.9775 0.7375 1.0475 0.7375 1.0475 0.635 1.1125 0.635 1.205 0.635 1.205 0.7 1.1125 0.7 1.1125 0.7375 1.1125 0.8025 0.9775 0.8025  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.85 0.54 2.4425 0.54 2.4425 0.675 2.3075 0.675 2.3075 0.605 1.85 0.605  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.9625 0.67 2.0225 0.67 2.0275 0.67 2.115 0.67 2.115 0.735 2.0275 0.735 2.0275 0.8375 1.9625 0.8375  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.395 0.15 0.53 0.15 0.53 0.375 1.15 0.375 1.15 0.15 1.285 0.15 1.285 0.375 1.73 0.375 1.73 0.15 1.795 0.15 1.795 0.41 2.485 0.41 2.485 0.15 2.55 0.15 2.55 0.475 1.785 0.475 1.785 0.94 2.095 0.94 2.16 0.94 2.475 0.94 2.475 0.76 2.54 0.76 2.54 1.035 2.475 1.035 2.475 1.005 2.16 1.005 2.16 1.075 2.095 1.075 2.095 1.005 1.785 1.005 1.785 1.035 1.72 1.035 1.72 0.44 0.465 0.44 0.465 0.355 0.395 0.355  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.42 0.4 0.42 0.4 0.5225 0.4 0.555 0.335 0.555 0.335 0.5225 0.2175 0.5225  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.66 -0.085 2.66 0.085 2.205 0.085 2.205 0.345 2.07 0.345 2.07 0.085 1.665 0.085 1.665 0.31 1.53 0.31 1.53 0.085 0.905 0.085 0.905 0.31 0.77 0.31 0.77 0.085 0.115 0.085 0.115 0.345 0.05 0.345 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.91 0.505 1.485 0.505 1.485 0.64 1.4575 0.64 1.4575 0.6975 1.3925 0.6975 1.3925 0.57 0.975 0.57 0.975 0.64 0.91 0.64  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.5625 0.15 0.5625 0.15 0.5975 0.25 0.5975 0.25 0.6325 0.695 0.6325 0.695 0.5625 0.76 0.5625 0.76 0.6975 0.15 0.6975 0.0625 0.6975  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.765 0.87 0.765 0.87 0.905 1.565 0.905 1.565 0.765 1.63 0.765 1.63 1.04 1.565 1.04 1.565 0.97 0.87 0.97 0.87 1.165 1.285 1.165 1.285 1.23 0.805 1.23 0.805 0.83 0.485 0.83 0.485 1.04 0.42 1.04 0.42 0.83 0.11 0.83 0.11 1.04 0.045 1.04  ;
        POLYGON 0.955 1.035 1.09 1.035 1.375 1.035 1.44 1.035 1.44 1.1 1.44 1.14 1.905 1.14 1.905 1.07 1.97 1.07 1.97 1.14 2.285 1.14 2.285 1.07 2.35 1.07 2.35 1.205 2.285 1.205 1.97 1.205 1.905 1.205 1.375 1.205 1.375 1.1 1.09 1.1 0.955 1.1  ;
  END
END AOI222_X4

MACRO AOI22_X1
  CLASS core ;
  FOREIGN AOI22_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 1.0325 0.295 1.0325 0.295 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.7025 0.34 0.7025 0.34 0.8375 0.2525 0.8375  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.57 0.2825 0.6975 0.2825 0.6975 0.4975 0.57 0.4975  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.865 0.085 0.865 0.3175 0.8 0.3175 0.8 0.085 0.11 0.085 0.11 0.3175 0.045 0.3175 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.4225 0.1275 0.4225 0.1275 0.5575 0.0625 0.5575  ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.5625 0.785 0.5625 0.785 0.6975 0.6325 0.6975  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.425 0.2375 0.49 0.2375 0.49 0.5625 0.5075 0.5625 0.5075 0.7625 0.675 0.7625 0.675 1.045 0.61 1.045 0.61 0.8275 0.4575 0.8275 0.4575 0.805 0.425 0.805  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.9025 0.485 0.9025 0.485 1.11 0.8 1.11 0.8 1.0325 0.865 1.0325 0.865 1.175 0.42 1.175 0.42 0.9675 0.11 0.9675 0.11 1.045 0.045 1.045  ;
  END
END AOI22_X1

MACRO AOI22_X2
  CLASS core ;
  FOREIGN AOI22_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2525 1.315 0.2525 0.8925 0.3175 0.8925 0.3175 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.4225 0.3625 0.4225 0.3625 0.5575 0.2525 0.5575  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.5775 0.1775 0.7325 0.1775 0.7325 0.2425 0.6425 0.2425 0.6425 0.5575 0.5775 0.5575  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.8875 0.085 0.8875 0.3875 0.8225 0.3875 0.8225 0.085 0.1325 0.085 0.1325 0.3875 0.0675 0.3875 0.0675 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.5625 0.1275 0.5625 0.1275 0.6975 0.0625 0.6975  ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.7425 0.48 0.8075 0.48 0.8075 0.55 0.8875 0.55 0.8875 0.6975 0.8225 0.6975 0.8225 0.615 0.7425 0.615  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4475 0.1575 0.5125 0.1575 0.5125 0.6225 0.5975 0.6225 0.5975 0.645 0.6775 0.645 0.6775 0.6625 0.6975 0.6625 0.6975 0.9875 0.6325 0.9875 0.6325 0.71 0.5475 0.71 0.5475 0.6875 0.4475 0.6875  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.0675 0.7625 0.5075 0.7625 0.5075 1.0525 0.8225 1.0525 0.8225 0.8425 0.8875 0.8425 0.8875 1.1175 0.4425 1.1175 0.4425 0.8275 0.1325 0.8275 0.1325 1.0375 0.0675 1.0375  ;
  END
END AOI22_X2

MACRO AOI22_X4
  CLASS core ;
  FOREIGN AOI22_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.71 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2425 1.315 0.2425 1.025 0.3075 1.025 0.3075 1.315 0.6225 1.315 0.6225 1.025 0.6875 1.025 0.6875 1.315 1.71 1.315 1.71 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.4225 0.3625 0.4225 0.3625 0.5575 0.2525 0.5575  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.3475 0.2825 1.4575 0.2825 1.4575 0.4175 1.4125 0.4175 1.4125 0.55 1.3475 0.55  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.71 -0.085 1.71 0.085 1.6475 0.085 1.6475 0.38 1.5825 0.38 1.5825 0.085 0.8875 0.085 0.8875 0.38 0.8225 0.38 0.8225 0.085 0.1325 0.085 0.1325 0.38 0.0675 0.38 0.0675 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.5625 0.1275 0.5625 0.1275 0.6225 0.7775 0.6225 0.7775 0.7575 0.7125 0.7575 0.7125 0.6875 0.2275 0.6875 0.2275 0.7575 0.1625 0.7575 0.1625 0.6975 0.0625 0.6975  ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.9725 0.575 1.0375 0.575 1.0375 0.6325 1.4775 0.6325 1.4775 0.5625 1.6475 0.5625 1.6475 0.6975 1.0375 0.6975 1.0375 0.71 0.9725 0.71  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.9075 0.775 1.0775 0.775 1.0775 0.845 1.4575 0.845 1.4575 1.12 1.3925 1.12 1.3925 0.91 1.0775 0.91 1.0775 1.12 1.0125 1.12 1.0125 0.84 0.8425 0.84 0.8425 0.51 0.4475 0.51 0.4475 0.15 0.5125 0.15 0.5125 0.445 1.2025 0.445 1.2025 0.15 1.2675 0.15 1.2675 0.51 0.9075 0.51  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.0575 0.895 0.8075 0.895 0.8075 0.935 0.8775 0.935 0.8775 1.185 1.2025 1.185 1.2025 0.975 1.2675 0.975 1.2675 1.185 1.5825 1.185 1.5825 0.975 1.6475 0.975 1.6475 1.25 0.8125 1.25 0.8125 1 0.7475 1 0.7475 0.96 0.4975 0.96 0.4975 1.17 0.4325 1.17 0.4325 0.96 0.1225 0.96 0.1225 1.17 0.0575 1.17  ;
  END
END AOI22_X4

MACRO BUF_X1
  CLASS core ;
  FOREIGN BUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.7375 0.42 0.7375 0.42 0.1525 0.485 0.1525 0.485 0.9425 0.42 0.9425 0.42 0.8025 0.2175 0.8025  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.5375 0.24 0.5375 0.24 0.5975 0.3525 0.5975 0.3525 0.6625 0.24 0.6625 0.24 0.6725 0.175 0.6725  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 0.8675 0.295 0.8675 0.295 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.295 0.085 0.295 0.2725 0.23 0.2725 0.23 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.1525 0.11 0.1525 0.11 0.4075 0.29 0.4075 0.29 0.3375 0.355 0.3375 0.355 0.4725 0.11 0.4725 0.11 0.9425 0.045 0.9425  ;
  END
END BUF_X1

MACRO BUF_X16
  CLASS core ;
  FOREIGN BUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.53 0.5975 0.905 0.5975 0.905 0.9875 0.84 0.9875 0.84 0.6625 0.53 0.6625 0.53 0.9875 0.465 0.9875 0.465 0.2025 0.53 0.2025 0.53 0.3975 0.84 0.3975 0.84 0.1875 0.905 0.1875 0.905 0.4625 0.53 0.4625  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2 0.5875 0.265 0.5875 0.265 0.7375 0.3525 0.7375 0.3525 0.8025 0.2 0.8025  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.275 1.315 0.275 1.0375 0.34 1.0375 0.34 1.315 0.65 1.315 0.65 1.0375 0.715 1.0375 0.715 1.315 1.03 1.315 1.03 1.0375 1.095 1.0375 1.095 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 1.095 0.085 1.095 0.3325 1.03 0.3325 1.03 0.085 0.715 0.085 0.715 0.3325 0.65 0.3325 0.65 0.085 0.34 0.085 0.34 0.3325 0.275 0.3325 0.275 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.07 0.3425 0.135 0.3425 0.135 0.4575 0.4 0.4575 0.4 0.6025 0.335 0.6025 0.335 0.5225 0.135 0.5225 0.135 0.8475 0.07 0.8475  ;
  END
END BUF_X16

MACRO BUF_X2
  CLASS core ;
  FOREIGN BUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.7375 0.435 0.7375 0.435 0.2125 0.5 0.2125 0.5 1.0875 0.435 1.0875 0.435 0.8025 0.2175 0.8025  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.5375 0.24 0.5375 0.24 0.5975 0.3525 0.5975 0.3525 0.6625 0.24 0.6625 0.24 0.6725 0.175 0.6725  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.25 1.315 0.25 0.8675 0.315 0.8675 0.315 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.31 0.085 0.31 0.2725 0.245 0.2725 0.245 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.43 0.06 0.43 0.06 0.1525 0.125 0.1525 0.125 0.4075 0.305 0.4075 0.305 0.3375 0.37 0.3375 0.37 0.4725 0.11 0.4725 0.11 1.0825 0.045 1.0825  ;
  END
END BUF_X2

MACRO BUF_X32
  CLASS core ;
  FOREIGN BUF_X32 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.71 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.53 0.7375 1.665 0.7375 1.665 1.0125 1.6 1.0125 1.6 0.8025 1.285 0.8025 1.285 1.0125 1.22 1.0125 1.22 0.8025 0.905 0.8025 0.905 1.0125 0.84 1.0125 0.84 0.8025 0.53 0.8025 0.53 0.94 0.465 0.94 0.465 0.2675 0.53 0.2675 0.53 0.41 0.84 0.41 0.84 0.2 0.905 0.2 0.905 0.41 1.22 0.41 1.22 0.2 1.285 0.2 1.285 0.41 1.6 0.41 1.6 0.2 1.665 0.2 1.665 0.475 0.53 0.475  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.185 0.54 0.25 0.54 0.25 0.7375 0.3525 0.7375 0.3525 0.8025 0.185 0.8025  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.275 1.315 0.275 1.0675 0.34 1.0675 0.34 1.315 0.65 1.315 0.65 1.0675 0.715 1.0675 0.715 1.315 1.03 1.315 1.03 1.0675 1.095 1.0675 1.095 1.315 1.41 1.315 1.41 1.0675 1.475 1.0675 1.475 1.315 1.71 1.315 1.71 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.71 -0.085 1.71 0.085 1.475 0.085 1.475 0.345 1.41 0.345 1.41 0.085 1.095 0.085 1.095 0.345 1.03 0.345 1.03 0.085 0.715 0.085 0.715 0.345 0.65 0.345 0.65 0.085 0.34 0.085 0.34 0.345 0.275 0.345 0.275 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.055 0.4325 0.07 0.4325 0.07 0.21 0.135 0.21 0.135 0.41 0.375 0.41 0.375 0.4225 0.4 0.4225 0.4 0.6675 0.335 0.6675 0.335 0.475 0.12 0.475 0.12 0.8 0.055 0.8  ;
  END
END BUF_X32

MACRO BUF_X4
  CLASS core ;
  FOREIGN BUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.8775 0.435 0.8775 0.435 0.225 0.5 0.225 0.5 1.0175 0.435 1.0175 0.435 0.9425 0.2175 0.9425  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.6175 0.24 0.6175 0.24 0.7375 0.3525 0.7375 0.3525 0.8025 0.175 0.8025  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.25 1.315 0.25 1.0675 0.315 1.0675 0.315 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.315 0.085 0.315 0.355 0.25 0.355 0.25 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.365 0.11 0.365 0.11 0.4875 0.37 0.4875 0.37 0.625 0.305 0.625 0.305 0.5525 0.11 0.5525 0.11 0.8775 0.045 0.8775  ;
  END
END BUF_X4

MACRO BUF_X8
  CLASS core ;
  FOREIGN BUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.225 0.5075 0.225 0.5075 1.0175 0.4425 1.0175  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1825 0.6175 0.2475 0.6175 0.2475 0.8425 0.3175 0.8425 0.3175 0.9775 0.1825 0.9775  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2575 1.315 0.2575 1.0675 0.3225 1.0675 0.3225 1.315 0.6325 1.315 0.6325 1.0675 0.6975 1.0675 0.6975 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.6975 0.085 0.6975 0.355 0.6325 0.355 0.6325 0.085 0.3225 0.085 0.3225 0.355 0.2575 0.355 0.2575 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.0525 0.365 0.1175 0.365 0.1175 0.4875 0.3775 0.4875 0.3775 0.625 0.3125 0.625 0.3125 0.5525 0.1175 0.5525 0.1175 0.8775 0.0525 0.8775  ;
  END
END BUF_X8

MACRO CLKBUF_X1
  CLASS core ;
  FOREIGN CLKBUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.7375 0.42 0.7375 0.42 0.1525 0.485 0.1525 0.485 0.9425 0.42 0.9425 0.42 0.8025 0.2175 0.8025  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.5375 0.24 0.5375 0.24 0.5975 0.3525 0.5975 0.3525 0.6625 0.24 0.6625 0.24 0.6725 0.175 0.6725  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 0.8675 0.295 0.8675 0.295 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.295 0.085 0.295 0.2725 0.23 0.2725 0.23 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.1525 0.11 0.1525 0.11 0.4075 0.29 0.4075 0.29 0.3375 0.355 0.3375 0.355 0.4725 0.11 0.4725 0.11 0.9425 0.045 0.9425  ;
  END
END CLKBUF_X1

MACRO CLKBUF_X2
  CLASS core ;
  FOREIGN CLKBUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.7375 0.435 0.7375 0.435 0.2125 0.5 0.2125 0.5 1.0875 0.435 1.0875 0.435 0.8025 0.2175 0.8025  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.5375 0.24 0.5375 0.24 0.5975 0.3525 0.5975 0.3525 0.6625 0.24 0.6625 0.24 0.6725 0.175 0.6725  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.25 1.315 0.25 0.8675 0.315 0.8675 0.315 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.31 0.085 0.31 0.2725 0.245 0.2725 0.245 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.43 0.06 0.43 0.06 0.1525 0.125 0.1525 0.125 0.4075 0.305 0.4075 0.305 0.3375 0.37 0.3375 0.37 0.4725 0.11 0.4725 0.11 1.0825 0.045 1.0825  ;
  END
END CLKBUF_X2

MACRO CLKBUF_X3
  CLASS core ;
  FOREIGN CLKBUF_X3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.235 0.5075 0.235 0.5075 1.12 0.4425 1.12  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1825 0.72 0.2475 0.72 0.2475 0.8775 0.3525 0.8775 0.3525 0.9425 0.1825 0.9425  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2575 1.315 0.2575 1.035 0.3225 1.035 0.3225 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.3225 0.085 0.3225 0.455 0.2575 0.455 0.2575 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.0525 0.375 0.1175 0.375 0.1175 0.59 0.3125 0.59 0.3125 0.52 0.3775 0.52 0.3775 0.655 0.1175 0.655 0.1175 1.25 0.0525 1.25  ;
  END
END CLKBUF_X3

MACRO CLKGATETST_X1
  CLASS core ;
  FOREIGN CLKGATETST_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.85 BY 1.4 ;
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.4 0.105 0.4 0.105 0.3375 0.17 0.3375 0.17 0.4725 0.1275 0.4725 0.1275 0.5575 0.0625 0.5575  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.42 1.315 0.42 0.9425 0.485 0.9425 0.485 1.315 1.18 1.315 1.18 0.9425 1.245 0.9425 1.245 1.315 1.73 1.315 1.73 0.845 1.795 0.845 1.795 1.315 2.075 1.315 2.075 0.9025 2.14 0.9025 2.14 1.315 2.45 1.315 2.45 0.9025 2.515 0.9025 2.515 1.315 2.85 1.315 2.85 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.85 -0.085 2.85 0.085 2.55 0.085 2.55 0.375 2.415 0.375 2.415 0.085 1.795 0.085 1.795 0.445 1.73 0.445 1.73 0.085 1.245 0.085 1.245 0.2425 1.18 0.2425 1.18 0.085 0.485 0.085 0.485 0.2425 0.42 0.2425 0.42 0.085 0.11 0.085 0.11 0.2425 0.045 0.2425 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN GCK
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.5325 0.7025 2.64 0.7025 2.64 0.29 2.72 0.29 2.72 1.1625 2.655 1.1625 2.655 0.8375 2.5325 0.8375  ;
    END
  END GCK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3575 0.6675 0.445 0.6675 0.445 0.7025 0.5075 0.7025 0.5075 0.8375 0.3575 0.8375  ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.1175 0.5975 2.2525 0.5975 2.2525 0.6625 2.2 0.6625 2.2 0.7675 2.1175 0.7675  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.7575 0.2275 0.7575 0.2275 0.57 0.235 0.57 0.235 0.2125 0.3 0.2125 0.3 0.4075 0.5 0.4075 0.5 0.3375 0.565 0.3375 0.565 0.4725 0.3 0.4725 0.3 0.6025 0.2925 0.6025 0.2925 0.8225 0.11 0.8225 0.11 1.0675 0.045 1.0675  ;
        POLYGON 0.695 0.8125 1.24 0.8125 1.24 0.7425 1.305 0.7425 1.305 0.8775 0.865 0.8775 0.865 1.1625 0.8 1.1625 0.8 0.9175 0.63 0.9175 0.63 0.1925 0.8 0.1925 0.8 0.155 0.865 0.155 0.865 0.29 0.695 0.29  ;
        POLYGON 1.1 0.4075 1.37 0.4075 1.37 0.2125 1.435 0.2125 1.435 0.4125 1.48 0.4125 1.48 0.5475 1.41 0.5475 1.41 0.4725 1.165 0.4725 1.165 0.5425 1.1 0.5425  ;
        POLYGON 1.37 0.7425 1.48 0.7425 1.48 0.8775 1.435 0.8775 1.435 1.1625 1.37 1.1625  ;
        POLYGON 0.76 0.6125 0.91 0.6125 0.91 0.3375 0.975 0.3375 0.975 0.6125 1.545 0.6125 1.545 0.31 1.61 0.31 1.61 1.12 1.545 1.12 1.545 0.6775 0.825 0.6775 0.825 0.7475 0.76 0.7475  ;
        POLYGON 1.675 0.54 1.74 0.54 1.74 0.61 1.92 0.61 1.92 0.415 1.985 0.415 1.985 1.065 1.92 1.065 1.92 0.675 1.675 0.675  ;
        POLYGON 2.265 0.7675 2.385 0.7675 2.385 0.5325 2.075 0.5325 2.075 0.38 2.14 0.38 2.14 0.4675 2.575 0.4675 2.575 0.6375 2.45 0.6375 2.45 0.8325 2.33 0.8325 2.33 1.1225 2.265 1.1225  ;
  END
END CLKGATETST_X1

MACRO CLKGATETST_X2
  CLASS core ;
  FOREIGN CLKGATETST_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.85 BY 1.4 ;
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.4 0.105 0.4 0.105 0.3375 0.17 0.3375 0.17 0.4725 0.1275 0.4725 0.1275 0.5575 0.0625 0.5575  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.42 1.315 0.42 0.9425 0.485 0.9425 0.485 1.315 1.18 1.315 1.18 0.9425 1.245 0.9425 1.245 1.315 1.73 1.315 1.73 0.845 1.795 0.845 1.795 1.315 2.075 1.315 2.075 0.9025 2.14 0.9025 2.14 1.315 2.45 1.315 2.45 0.9025 2.515 0.9025 2.515 1.315 2.85 1.315 2.85 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.85 -0.085 2.85 0.085 2.55 0.085 2.55 0.375 2.415 0.375 2.415 0.085 1.795 0.085 1.795 0.445 1.73 0.445 1.73 0.085 1.245 0.085 1.245 0.2425 1.18 0.2425 1.18 0.085 0.485 0.085 0.485 0.2425 0.42 0.2425 0.42 0.085 0.11 0.085 0.11 0.2425 0.045 0.2425 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN GCK
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.655 1.0275 2.7225 1.0275 2.7225 0.8375 2.5325 0.8375 2.5325 0.7025 2.7225 0.7025 2.7225 0.425 2.64 0.425 2.64 0.36 2.64 0.29 2.72 0.29 2.72 0.36 2.7875 0.36 2.7875 0.425 2.7875 1.0275 2.7875 1.0925 2.72 1.0925 2.72 1.1625 2.655 1.1625 2.655 1.0925  ;
    END
  END GCK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3575 0.6675 0.445 0.6675 0.445 0.7025 0.5075 0.7025 0.5075 0.8375 0.3575 0.8375  ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.1175 0.5975 2.2525 0.5975 2.2525 0.6625 2.2 0.6625 2.2 0.7675 2.1175 0.7675  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.7575 0.2275 0.7575 0.2275 0.57 0.235 0.57 0.235 0.2125 0.3 0.2125 0.3 0.4075 0.5 0.4075 0.5 0.3375 0.565 0.3375 0.565 0.4725 0.3 0.4725 0.3 0.6025 0.2925 0.6025 0.2925 0.8225 0.11 0.8225 0.11 1.0675 0.045 1.0675  ;
        POLYGON 0.695 0.8125 1.24 0.8125 1.24 0.7425 1.305 0.7425 1.305 0.8775 0.865 0.8775 0.865 1.1625 0.8 1.1625 0.8 0.9175 0.63 0.9175 0.63 0.1925 0.8 0.1925 0.8 0.155 0.865 0.155 0.865 0.29 0.695 0.29  ;
        POLYGON 1.1 0.4075 1.37 0.4075 1.37 0.2125 1.435 0.2125 1.435 0.4125 1.48 0.4125 1.48 0.5475 1.41 0.5475 1.41 0.4725 1.165 0.4725 1.165 0.5425 1.1 0.5425  ;
        POLYGON 1.37 0.7425 1.48 0.7425 1.48 0.8775 1.435 0.8775 1.435 1.1625 1.37 1.1625  ;
        POLYGON 0.76 0.6125 0.91 0.6125 0.91 0.3375 0.975 0.3375 0.975 0.6125 1.545 0.6125 1.545 0.31 1.61 0.31 1.61 1.12 1.545 1.12 1.545 0.6775 0.825 0.6775 0.825 0.7475 0.76 0.7475  ;
        POLYGON 1.675 0.54 1.74 0.54 1.74 0.61 1.92 0.61 1.92 0.415 1.985 0.415 1.985 1.065 1.92 1.065 1.92 0.675 1.675 0.675  ;
        POLYGON 2.265 0.7675 2.385 0.7675 2.385 0.5325 2.075 0.5325 2.075 0.38 2.14 0.38 2.14 0.4675 2.45 0.4675 2.45 0.57 2.61 0.57 2.61 0.635 2.45 0.635 2.45 0.8325 2.33 0.8325 2.33 1.1225 2.265 1.1225  ;
  END
END CLKGATETST_X2

MACRO CLKGATETST_X4
  CLASS core ;
  FOREIGN CLKGATETST_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.85 BY 1.4 ;
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.4 0.105 0.4 0.105 0.3375 0.17 0.3375 0.17 0.4725 0.1275 0.4725 0.1275 0.5575 0.0625 0.5575  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.42 1.315 0.42 0.9425 0.485 0.9425 0.485 1.315 1.18 1.315 1.18 0.9425 1.245 0.9425 1.245 1.315 1.73 1.315 1.73 0.845 1.795 0.845 1.795 1.315 2.075 1.315 2.075 0.99 2.14 0.99 2.14 1.315 2.45 1.315 2.45 0.99 2.515 0.99 2.515 1.315 2.85 1.315 2.85 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.85 -0.085 2.85 0.085 2.55 0.085 2.55 0.375 2.415 0.375 2.415 0.085 1.795 0.085 1.795 0.445 1.73 0.445 1.73 0.085 1.245 0.085 1.245 0.2425 1.18 0.2425 1.18 0.085 0.485 0.085 0.485 0.2425 0.42 0.2425 0.42 0.085 0.11 0.085 0.11 0.2425 0.045 0.2425 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN GCK
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.5325 0.7025 2.675 0.7025 2.675 0.4325 2.64 0.4325 2.64 0.1575 2.705 0.1575 2.705 0.3675 2.74 0.3675 2.74 0.7675 2.705 0.7675 2.705 0.86 2.705 0.8625 2.705 1.1225 2.64 1.1225 2.64 0.8625 2.64 0.86 2.64 0.8375 2.5325 0.8375  ;
    END
  END GCK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3575 0.6675 0.445 0.6675 0.445 0.7025 0.5075 0.7025 0.5075 0.8375 0.3575 0.8375  ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.1175 0.5975 2.2525 0.5975 2.2525 0.6625 2.2 0.6625 2.2 0.7675 2.1175 0.7675  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.7575 0.2275 0.7575 0.2275 0.57 0.235 0.57 0.235 0.2125 0.3 0.2125 0.3 0.4075 0.5 0.4075 0.5 0.3375 0.565 0.3375 0.565 0.4725 0.3 0.4725 0.3 0.6025 0.2925 0.6025 0.2925 0.8225 0.11 0.8225 0.11 1.0675 0.045 1.0675  ;
        POLYGON 0.695 0.8125 1.24 0.8125 1.24 0.7425 1.305 0.7425 1.305 0.8775 0.865 0.8775 0.865 1.1625 0.8 1.1625 0.8 0.9175 0.63 0.9175 0.63 0.1925 0.8 0.1925 0.8 0.155 0.865 0.155 0.865 0.29 0.695 0.29  ;
        POLYGON 1.1 0.4075 1.37 0.4075 1.37 0.2125 1.435 0.2125 1.435 0.4125 1.48 0.4125 1.48 0.5475 1.41 0.5475 1.41 0.4725 1.165 0.4725 1.165 0.5425 1.1 0.5425  ;
        POLYGON 1.37 0.7425 1.48 0.7425 1.48 0.8775 1.435 0.8775 1.435 1.1625 1.37 1.1625  ;
        POLYGON 0.76 0.6125 0.91 0.6125 0.91 0.3375 0.975 0.3375 0.975 0.6125 1.545 0.6125 1.545 0.31 1.61 0.31 1.61 1.12 1.545 1.12 1.545 0.6775 0.825 0.6775 0.825 0.7475 0.76 0.7475  ;
        POLYGON 1.675 0.54 1.74 0.54 1.74 0.61 1.92 0.61 1.92 0.415 1.985 0.415 1.985 1.065 1.92 1.065 1.92 0.675 1.675 0.675  ;
        POLYGON 2.265 0.7675 2.385 0.7675 2.385 0.5325 2.075 0.5325 2.075 0.24 2.14 0.24 2.14 0.4675 2.45 0.4675 2.45 0.5725 2.61 0.5725 2.61 0.6375 2.45 0.6375 2.45 0.8325 2.33 0.8325 2.33 0.86 2.33 0.8625 2.33 1.1225 2.265 1.1225 2.265 0.8625 2.265 0.86  ;
  END
END CLKGATETST_X4

MACRO CLKGATETST_X8
  CLASS core ;
  FOREIGN CLKGATETST_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.04 BY 1.4 ;
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.4225 0.1275 0.4225 0.1275 0.5575 0.0625 0.5575  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.42 1.315 0.42 1.1575 0.485 1.1575 0.485 1.315 1.18 1.315 1.18 1.0175 1.245 1.0175 1.245 1.315 1.725 1.315 1.725 0.9025 1.79 0.9025 1.79 1.315 2.07 1.315 2.07 0.7 2.135 0.7 2.135 1.315 2.495 1.315 2.495 0.745 2.58 0.745 2.58 1.315 2.9025 1.315 2.9025 1.025 2.9675 1.025 2.9675 1.315 3.04 1.315 3.04 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.04 -0.085 3.04 0.085 2.99 0.085 2.99 0.3325 2.925 0.3325 2.925 0.085 2.58 0.085 2.58 0.4325 2.515 0.4325 2.515 0.085 1.795 0.085 1.795 0.34 1.73 0.34 1.73 0.085 1.245 0.085 1.245 0.3175 1.18 0.3175 1.18 0.085 0.485 0.085 0.485 0.3175 0.42 0.3175 0.42 0.085 0.11 0.085 0.11 0.3175 0.045 0.3175 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN GCK
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.7175 0.6725 2.7225 0.6725 2.7225 0.2025 2.8 0.2025 2.8 0.6975 2.7825 0.6975 2.7825 1.155 2.7175 1.155  ;
    END
  END GCK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3575 0.6125 0.4225 0.6125 0.4225 0.6825 0.5075 0.6825 0.5075 0.8375 0.4425 0.8375 0.4425 0.7475 0.3575 0.7475  ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.7725 0.4225 1.84 0.4225 1.84 0.57 1.7725 0.57  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.6525 0.055 0.6525 0.055 0.6225 0.2275 0.6225 0.2275 0.5275 0.23 0.5275 0.23 0.2875 0.295 0.2875 0.295 0.4825 0.5 0.4825 0.5 0.4125 0.565 0.4125 0.565 0.5475 0.2925 0.5475 0.2925 0.6875 0.11 0.6875 0.11 1.0125 0.045 1.0125  ;
        POLYGON 0.695 0.8875 0.8 0.8875 1.24 0.8875 1.24 0.8175 1.305 0.8175 1.305 0.9525 0.865 0.9525 0.865 1.2375 0.8 1.2375 0.8 0.9925 0.63 0.9925 0.63 0.8875 0.63 0.365 0.63 0.2675 0.8 0.2675 0.8 0.23 0.865 0.23 0.865 0.365 0.8 0.365 0.695 0.365  ;
        POLYGON 1.1 0.4125 1.37 0.4125 1.37 0.2725 1.435 0.2725 1.435 0.4125 1.48 0.4125 1.48 0.5475 1.415 0.5475 1.415 0.4775 1.165 0.4775 1.165 0.5475 1.1 0.5475  ;
        POLYGON 1.37 0.7425 1.48 0.7425 1.48 0.8775 1.435 0.8775 1.435 1.2375 1.37 1.2375  ;
        POLYGON 1.54 0.9025 1.545 0.9025 1.545 0.6775 0.825 0.6775 0.825 0.8225 0.76 0.8225 0.76 0.6125 0.91 0.6125 0.91 0.4125 0.975 0.4125 0.975 0.6125 1.545 0.6125 1.545 0.31 1.61 0.31 1.61 1.1775 1.54 1.1775  ;
        POLYGON 1.675 0.6275 1.74 0.6275 1.74 0.6975 1.92 0.6975 1.92 0.31 1.985 0.31 1.985 0.7225 1.98 0.7225 1.98 1.1225 1.915 1.1225 1.915 0.7625 1.675 0.7625  ;
        POLYGON 2.1 0.15 2.165 0.15 2.165 0.53 2.35 0.53 2.35 0.57 2.5925 0.57 2.5925 0.5 2.6575 0.5 2.6575 0.635 2.355 0.635 2.355 1.21 2.29 1.21 2.29 0.595 2.11 0.595 2.11 0.565 2.1 0.565  ;
  END
END CLKGATETST_X8

MACRO CLKGATE_X1
  CLASS core ;
  FOREIGN CLKGATE_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.47 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 0.8125 0.295 0.8125 0.295 1.315 0.99 1.315 0.99 0.8125 1.055 0.8125 1.055 1.315 1.675 1.315 1.675 0.8975 1.74 0.8975 1.74 1.315 2.05 1.315 2.05 0.8975 2.115 0.8975 2.115 1.315 2.18 1.315 2.47 1.315 2.47 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.47 -0.085 2.47 0.085 2.115 0.085 2.115 0.2975 2.05 0.2975 2.05 0.085 1.585 0.085 1.585 0.4475 1.52 0.4475 1.52 0.085 1.055 0.085 1.055 0.3175 0.99 0.3175 0.99 0.085 0.295 0.085 0.295 0.3175 0.23 0.3175 0.23 0.085 0 0.085  ;
    END
  END VSS
  PIN GCK
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.1525 0.5625 2.24 0.5625 2.24 0.1775 2.32 0.1775 2.32 1.1575 2.255 1.1575 2.255 0.6975 2.1525 0.6975  ;
    END
  END GCK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.8225 0.4225 0.91 0.4225 0.91 0.5575 0.8225 0.5575  ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.565 0.7025 1.6475 0.7025 1.6475 0.8375 1.565 0.8375  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.2875 0.11 0.2875 0.11 0.4825 0.315 0.4825 0.315 0.4125 0.38 0.4125 0.38 0.5475 0.11 0.5475 0.11 1.0325 0.045 1.0325  ;
        POLYGON 0.175 0.6125 0.24 0.6125 0.24 0.6825 0.61 0.6825 0.61 0.2875 0.675 0.2875 0.675 1.0325 0.61 1.0325 0.61 0.7475 0.175 0.7475  ;
        POLYGON 0.74 0.6225 1.18 0.6225 1.18 0.2875 1.245 0.2875 1.245 1.0325 1.18 1.0325 1.18 0.6875 0.805 0.6875 0.805 0.7575 0.74 0.7575  ;
        POLYGON 1.335 0.4175 1.4 0.4175 1.4 0.9025 1.55 0.9025 1.55 1.0375 1.485 1.0375 1.485 0.9675 1.335 0.9675  ;
        POLYGON 1.675 0.24 1.74 0.24 1.74 0.3325 1.925 0.3325 1.925 0.4325 2.11 0.4325 2.11 0.3625 2.175 0.3625 2.175 0.4975 1.925 0.4975 1.925 1.1175 1.86 1.1175 1.86 0.3975 1.69 0.3975 1.69 0.375 1.675 0.375  ;
  END
END CLKGATE_X1

MACRO CLKGATE_X2
  CLASS core ;
  FOREIGN CLKGATE_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.47 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 0.8125 0.295 0.8125 0.295 1.315 0.99 1.315 0.99 0.8125 1.055 0.8125 1.055 1.315 1.675 1.315 1.675 0.8975 1.74 0.8975 1.74 1.315 2.05 1.315 2.05 0.8975 2.115 0.8975 2.115 1.315 2.18 1.315 2.47 1.315 2.47 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.47 -0.085 2.47 0.085 2.115 0.085 2.115 0.2675 2.05 0.2675 2.05 0.085 1.585 0.085 1.585 0.1925 1.52 0.1925 1.52 0.085 1.055 0.085 1.055 0.3175 0.99 0.3175 0.99 0.085 0.295 0.085 0.295 0.3175 0.23 0.3175 0.23 0.085 0 0.085  ;
    END
  END VSS
  PIN GCK
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.1525 0.5625 2.24 0.5625 2.24 0.2375 2.32 0.2375 2.32 1.0675 2.255 1.0675 2.255 0.6975 2.1525 0.6975  ;
    END
  END GCK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.8225 0.4225 0.91 0.4225 0.91 0.5575 0.8225 0.5575  ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.565 0.7025 1.6475 0.7025 1.6475 0.8375 1.565 0.8375  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.2875 0.11 0.2875 0.11 0.4825 0.315 0.4825 0.315 0.4125 0.38 0.4125 0.38 0.5475 0.11 0.5475 0.11 1.0325 0.045 1.0325  ;
        POLYGON 0.175 0.6125 0.24 0.6125 0.24 0.6825 0.61 0.6825 0.61 0.2875 0.675 0.2875 0.675 1.0325 0.61 1.0325 0.61 0.7475 0.175 0.7475  ;
        POLYGON 0.74 0.6225 1.18 0.6225 1.18 0.2875 1.245 0.2875 1.245 1.0325 1.18 1.0325 1.18 0.6875 0.805 0.6875 0.805 0.7575 0.74 0.7575  ;
        POLYGON 1.335 0.1625 1.4 0.1625 1.4 0.9025 1.55 0.9025 1.55 1.0375 1.485 1.0375 1.485 0.9675 1.335 0.9675  ;
        POLYGON 1.675 0.2375 1.74 0.2375 1.74 0.33 1.925 0.33 1.925 0.4325 2.11 0.4325 2.11 0.3625 2.175 0.3625 2.175 0.4975 1.925 0.4975 1.925 1.1175 1.86 1.1175 1.86 0.395 1.69 0.395 1.69 0.3725 1.675 0.3725  ;
  END
END CLKGATE_X2

MACRO CLKGATE_X4
  CLASS core ;
  FOREIGN CLKGATE_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.47 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 0.8125 0.295 0.8125 0.295 1.315 0.99 1.315 0.99 0.8125 1.055 0.8125 1.055 1.315 1.6625 1.315 1.6625 0.9175 1.7275 0.9175 1.7275 1.315 2.015 1.315 2.015 0.9025 2.145 0.9025 2.15 0.9025 2.15 1.315 2.47 1.315 2.47 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.47 -0.085 2.47 0.085 2.135 0.085 2.135 0.3675 2.07 0.3675 2.07 0.085 1.585 0.085 1.585 0.1925 1.52 0.1925 1.52 0.085 1.055 0.085 1.055 0.3175 0.99 0.3175 0.99 0.085 0.295 0.085 0.295 0.3175 0.23 0.3175 0.23 0.085 0 0.085  ;
    END
  END VSS
  PIN GCK
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.1525 0.7025 2.255 0.7025 2.255 0.2375 2.32 0.2375 2.32 1.1375 2.255 1.1375 2.255 0.8375 2.1525 0.8375  ;
    END
  END GCK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.8225 0.4225 0.91 0.4225 0.91 0.5575 0.8225 0.5575  ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.5825 0.7025 1.6475 0.7025 1.6475 0.8375 1.5825 0.8375  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.2875 0.11 0.2875 0.11 0.4825 0.315 0.4825 0.315 0.4125 0.38 0.4125 0.38 0.5475 0.11 0.5475 0.11 1.0325 0.045 1.0325  ;
        POLYGON 0.175 0.6125 0.61 0.6125 0.61 0.2875 0.675 0.2875 0.675 1.0325 0.61 1.0325 0.61 0.6775 0.24 0.6775 0.24 0.7475 0.175 0.7475  ;
        POLYGON 0.74 0.6225 1.18 0.6225 1.18 0.2875 1.245 0.2875 1.245 1.0325 1.18 1.0325 1.18 0.6875 0.805 0.6875 0.805 0.7575 0.74 0.7575  ;
        POLYGON 1.335 0.1625 1.4 0.1625 1.4 0.49 1.5175 0.49 1.5175 1.1375 1.4525 1.1375 1.4525 0.555 1.335 0.555  ;
        POLYGON 1.675 0.1975 1.74 0.1975 1.74 0.5725 2.125 0.5725 2.125 0.5025 2.19 0.5025 2.19 0.6375 1.925 0.6375 1.925 1.1375 1.86 1.1375 1.86 0.6375 1.69 0.6375 1.69 0.615 1.675 0.615  ;
  END
END CLKGATE_X4

MACRO CLKGATE_X8
  CLASS core ;
  FOREIGN CLKGATE_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.66 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.7775 1.315 2.1175 1.315 2.1175 0.7275 2.2525 0.7275 2.2525 1.315 2.5375 1.315 2.5375 0.8325 2.6025 0.8325 2.6025 1.315 2.66 1.315 2.66 1.485 0 1.485 0 1.315 0.3225 1.315 0.3225 0.9025 0.2875 0.9025 0.2875 0.8375 0.4225 0.8375 0.4225 0.9025 0.3875 0.9025 0.3875 1.315 1.0825 1.315 1.0825 1.0425 1.0475 1.0425 1.0475 0.8375 1.1825 0.8375 1.1825 1.0425 1.1475 1.0425 1.1475 1.315 1.7125 1.315 1.7125 0.8425 1.6925 0.8425 1.6925 0.7775 1.8275 0.7775 1.8275 0.8425 1.7775 0.8425  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.0475 0.2625 1.1175 0.2625 1.1175 0.085 0.4225 0.085 0.4225 0.3275 0.2875 0.3275 0.2875 0.2625 0.3575 0.2625 0.3575 0.085 0 0.085 0 -0.085 2.66 -0.085 2.66 0.085 2.6025 0.085 2.6025 0.4075 2.5375 0.4075 2.5375 0.085 2.2625 0.085 2.2625 0.5125 2.1275 0.5125 2.1275 0.085 1.6775 0.085 1.6775 0.1525 1.6775 0.2325 1.6775 0.2675 1.6125 0.2675 1.6125 0.2325 1.6125 0.1525 1.6125 0.085 1.1825 0.085 1.1825 0.3275 1.0475 0.3275  ;
    END
  END VSS
  PIN GCK
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.3175 0.7225 2.3525 0.7225 2.3525 0.51 2.3525 0.4225 2.3425 0.4225 2.3425 0.2775 2.4175 0.2775 2.4175 0.4125 2.4175 0.4225 2.4175 0.51 2.4175 0.7225 2.4525 0.7225 2.4525 0.9275 2.3175 0.9275  ;
    END
  END GCK
  PIN E
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.9425 0.4925 1.0125 0.4925 1.0125 0.4225 1.0775 0.4225 1.0775 0.5575 0.9425 0.5575  ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.5775 0.4225 1.6475 0.4225 1.6475 0.4475 1.6725 0.4475 1.6725 0.5825 1.6475 0.5825 1.6075 0.5825 1.6075 0.5575 1.5775 0.5575  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.1375 0.3325 0.2025 0.3325 0.2025 0.4925 0.5075 0.4925 0.5075 0.5575 0.2025 0.5575 0.2025 1.0225 0.1375 1.0225  ;
        POLYGON 0.7325 0.7825 0.8025 0.7825 0.8025 0.9875 0.6675 0.9875 0.6675 0.7575 0.2825 0.7575 0.2825 0.6225 0.6675 0.6225 0.6675 0.3675 0.8025 0.3675 0.8025 0.4325 0.7325 0.4325  ;
        POLYGON 0.7975 0.6225 1.2725 0.6225 1.2725 0.3325 1.3375 0.3325 1.3375 1.0225 1.2725 1.0225 1.2725 0.6875 0.7975 0.6875  ;
        POLYGON 1.4275 0.2375 1.4925 0.2375 1.4925 0.35 1.4925 0.7225 1.6275 0.7225 1.6275 0.7875 1.4275 0.7875 1.4275 0.35  ;
        POLYGON 1.7675 0.2375 1.8325 0.2375 1.8325 0.5875 2.2875 0.5875 2.2875 0.6525 2.0275 0.6525 2.0275 0.9275 1.8925 0.9275 1.8925 0.6525 1.7675 0.6525  ;
  END
END CLKGATE_X8

MACRO DFFRS_X1
  CLASS core ;
  FOREIGN DFFRS_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 5.89 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 5.755 0.735 5.79 0.735 5.79 0.4175 5.755 0.4175 5.755 0.15 5.82 0.15 5.82 0.185 5.855 0.185 5.855 0.835 5.82 0.835 5.82 0.87 5.755 0.87  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.8 0.755 3.075 0.755 3.075 0.72 3.715 0.72 3.715 0.785 3.3925 0.785 3.3925 0.8025 3.2575 0.8025 3.2575 0.785 3.135 0.785 3.135 0.82 2.8 0.82  ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 4.01 0.75 4.455 0.75 4.455 0.955 4.39 0.955 4.39 0.815 3.945 0.815 3.945 0.65 3.91 0.65 3.91 0.585 3.945 0.585 3.945 0.425 3.645 0.425 3.645 0.27 2.885 0.27 2.885 0.425 2.49 0.425 2.49 0.27 2.095 0.27 2.095 0.59 1.75 0.59 1.75 0.525 2.03 0.525 2.03 0.205 2.1175 0.205 2.1175 0.1775 2.2525 0.1775 2.2525 0.205 2.555 0.205 2.555 0.36 2.82 0.36 2.82 0.205 3.71 0.205 3.71 0.36 4.01 0.36 4.01 0.585 4.045 0.585 4.045 0.65 4.01 0.65  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.42 1.315 4.13 1.315 4.13 1.06 4.195 1.06 4.195 1.315 4.85 1.315 4.85 0.685 4.95 0.685 4.95 1.315 5.23 1.315 5.23 0.685 5.295 0.685 5.295 1.315 5.57 1.315 5.57 0.795 5.635 0.795 5.635 1.315 5.89 1.315 5.89 1.485 0 1.485 0 1.315 0.275 1.315 0.275 0.9 0.34 0.9 0.34 1.315 1.03 1.315 1.03 1.155 1.095 1.155 1.095 1.315 1.89 1.315 1.89 1.075 1.955 1.075 1.955 1.315 2.635 1.315 2.635 1.13 2.6 1.13 2.6 1.065 2.735 1.065 2.735 1.13 2.7 1.13 2.7 1.315 3.355 1.315 3.355 1.175 3.32 1.175 3.32 1.11 3.455 1.11 3.455 1.175 3.42 1.175  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 5.3825 0.7025 5.415 0.7025 5.415 0.665 5.6 0.665 5.6 0.4 5.415 0.4 5.415 0.265 5.48 0.265 5.48 0.335 5.665 0.335 5.665 0.73 5.48 0.73 5.48 0.8 5.465 0.8 5.465 0.8375 5.3825 0.8375  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.775 0.23 3.81 0.23 3.81 0.085 2.72 0.085 2.72 0.23 2.755 0.23 2.755 0.295 2.62 0.295 2.62 0.23 2.655 0.23 2.655 0.085 1.93 0.085 1.93 0.35 1.965 0.35 1.965 0.415 1.83 0.415 1.83 0.35 1.865 0.35 1.865 0.085 0.7 0.085 0.7 0.26 0.735 0.26 0.735 0.325 0.635 0.325 0.6 0.325 0.6 0.26 0.635 0.26 0.635 0.085 0.34 0.085 0.34 0.235 0.34 0.39 0.275 0.39 0.275 0.235 0.275 0.085 0 0.085 0 -0.085 5.89 -0.085 5.89 0.085 5.635 0.085 5.635 0.27 5.57 0.27 5.57 0.085 5.295 0.085 5.295 0.4 5.23 0.4 5.23 0.085 3.875 0.085 3.875 0.23 3.91 0.23 3.91 0.295 3.775 0.295  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.4225 0.715 0.4225 0.715 0.68 0.6325 0.68  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.205 0.685 0.3525 0.685 0.3525 0.82 0.205 0.82  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.04 0.36 0.155 0.36 0.155 0.445 0.155 0.48 0.155 0.52 0.35 0.52 0.35 0.485 0.415 0.485 0.415 0.62 0.35 0.62 0.35 0.585 0.14 0.585 0.14 1.12 0.04 1.12 0.04 0.48 0.04 0.445  ;
        POLYGON 0.48 0.36 0.545 0.36 0.545 0.395 0.545 0.445 0.545 0.46 0.545 0.48 0.545 0.745 0.95 0.745 0.95 0.71 1.015 0.71 1.015 0.845 0.95 0.845 0.95 0.81 0.545 0.81 0.545 0.98 0.48 0.98 0.48 0.48 0.48 0.46 0.48 0.445 0.48 0.395  ;
        POLYGON 1.28 0.81 1.315 0.81 1.315 0.595 0.86 0.595 0.86 0.53 1.38 0.53 1.38 0.81 1.415 0.81 1.415 0.875 1.28 0.875  ;
        POLYGON 0.655 0.875 0.72 0.875 0.72 1.005 1.48 1.005 1.48 0.43 1.365 0.43 1.365 0.465 1.3 0.465 1.3 0.33 1.365 0.33 1.365 0.365 1.545 0.365 1.545 0.935 2.35 0.935 2.35 1.145 2.285 1.145 2.285 1 1.58 1 1.58 1.21 1.515 1.21 1.515 1.07 0.72 1.07 0.72 1.15 0.655 1.15  ;
        POLYGON 1.61 0.655 2.23 0.655 2.23 0.4 2.16 0.4 2.16 0.335 2.295 0.335 2.295 0.665 2.48 0.665 2.48 0.835 2.515 0.835 2.515 1.11 2.45 1.11 2.45 0.97 2.415 0.97 2.415 0.73 2.26 0.73 2.26 0.72 1.61 0.72  ;
        POLYGON 2.36 0.495 2.885 0.495 2.885 0.56 2.36 0.56  ;
        POLYGON 3.08 0.495 3.215 0.495 3.215 0.535 3.845 0.535 3.845 0.88 3.915 0.88 3.915 0.945 3.78 0.945 3.78 0.6 3.155 0.6 3.155 0.56 3.08 0.56  ;
        POLYGON 2.735 0.935 2.955 0.935 2.955 0.97 3.585 0.97 3.585 1.04 4 1.04 4 0.93 4.325 0.93 4.325 1.02 4.555 1.02 4.555 0.945 4.52 0.945 4.52 0.88 4.555 0.88 4.555 0.685 4.11 0.685 4.11 0.55 4.175 0.55 4.175 0.62 4.62 0.62 4.62 0.88 4.655 0.88 4.655 0.945 4.62 0.945 4.62 1.085 4.26 1.085 4.26 0.995 4.065 0.995 4.065 1.105 3.52 1.105 3.52 1.035 2.855 1.035 2.855 1 2.67 1 2.67 0.625 2.95 0.625 2.95 0.335 3.165 0.335 3.165 0.4 3.015 0.4 3.015 0.69 2.735 0.69  ;
        POLYGON 4.415 1.15 4.72 1.15 4.72 0.295 4.41 0.295 4.41 0.33 4.345 0.33 4.345 0.295 4.15 0.295 4.15 0.23 4.345 0.23 4.345 0.195 4.41 0.195 4.41 0.23 4.785 0.23 4.785 1.215 4.415 1.215  ;
        POLYGON 4.85 0.32 4.915 0.32 4.915 0.5 5.47 0.5 5.47 0.465 5.535 0.465 5.535 0.6 5.47 0.6 5.47 0.565 5.1 0.565 5.1 0.76 5.035 0.76 5.035 0.565 4.85 0.565  ;
  END
END DFFRS_X1

MACRO DFFRS_X2
  CLASS core ;
  FOREIGN DFFRS_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 5.89 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 5.7625 0.8425 5.7775 0.8425 5.7775 0.7425 5.7775 0.2675 5.7775 0.15 5.8425 0.15 5.8425 0.185 5.85 0.185 5.85 0.2675 5.85 0.7425 5.85 0.8425 5.85 0.9775 5.85 1.095 5.7775 1.095 5.7775 0.9775 5.7625 0.9775  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.8 0.755 3.075 0.755 3.075 0.72 3.715 0.72 3.715 0.785 3.3925 0.785 3.3925 0.8025 3.2575 0.8025 3.2575 0.785 3.135 0.785 3.135 0.82 2.8 0.82  ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 4.01 0.75 4.455 0.75 4.455 0.955 4.39 0.955 4.39 0.815 3.945 0.815 3.945 0.65 3.91 0.65 3.91 0.585 3.945 0.585 3.945 0.425 3.645 0.425 3.645 0.27 2.885 0.27 2.885 0.425 2.49 0.425 2.49 0.27 2.095 0.27 2.095 0.59 1.75 0.59 1.75 0.525 2.03 0.525 2.03 0.205 2.1175 0.205 2.1175 0.1775 2.2525 0.1775 2.2525 0.205 2.555 0.205 2.555 0.36 2.82 0.36 2.82 0.205 3.71 0.205 3.71 0.36 4.01 0.36 4.01 0.585 4.045 0.585 4.045 0.65 4.01 0.65  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.42 1.315 4.13 1.315 4.13 1.06 4.195 1.06 4.195 1.315 4.85 1.315 4.85 0.685 4.95 0.685 4.95 1.315 5.245 1.315 5.245 0.68 5.31 0.68 5.31 1.315 5.5925 1.315 5.5925 1.105 5.5925 0.94 5.5925 0.82 5.6575 0.82 5.6575 0.94 5.6575 1.105 5.6575 1.315 5.89 1.315 5.89 1.485 0 1.485 0 1.315 0.275 1.315 0.275 0.9 0.34 0.9 0.34 1.315 1.03 1.315 1.03 1.155 1.095 1.155 1.095 1.315 1.89 1.315 1.89 1.075 1.955 1.075 1.955 1.315 2.635 1.315 2.635 1.13 2.6 1.13 2.6 1.065 2.735 1.065 2.735 1.13 2.7 1.13 2.7 1.315 3.355 1.315 3.355 1.175 3.32 1.175 3.32 1.11 3.455 1.11 3.455 1.175 3.42 1.175  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 5.3825 0.7025 5.415 0.7025 5.415 0.665 5.43 0.665 5.58 0.665 5.6225 0.665 5.6225 0.4 5.58 0.4 5.515 0.4 5.5 0.4 5.43 0.4 5.43 0.265 5.495 0.265 5.495 0.335 5.5 0.335 5.515 0.335 5.58 0.335 5.6875 0.335 5.6875 0.73 5.58 0.73 5.5025 0.73 5.5025 0.94 5.43 0.94 5.43 0.8375 5.3825 0.8375  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.775 0.23 3.81 0.23 3.81 0.085 2.72 0.085 2.72 0.23 2.755 0.23 2.755 0.295 2.62 0.295 2.62 0.23 2.655 0.23 2.655 0.085 1.93 0.085 1.93 0.35 1.965 0.35 1.965 0.415 1.83 0.415 1.83 0.35 1.865 0.35 1.865 0.085 0.7 0.085 0.7 0.26 0.735 0.26 0.735 0.325 0.6 0.325 0.6 0.26 0.635 0.26 0.635 0.085 0.34 0.085 0.34 0.39 0.275 0.39 0.275 0.085 0 0.085 0 -0.085 5.89 -0.085 5.89 0.085 5.6575 0.085 5.6575 0.145 5.6575 0.27 5.5925 0.27 5.5925 0.145 5.5925 0.085 5.295 0.085 5.295 0.4 5.23 0.4 5.23 0.085 3.875 0.085 3.875 0.23 3.91 0.23 3.91 0.295 3.775 0.295  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.4225 0.715 0.4225 0.715 0.68 0.6325 0.68  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.205 0.685 0.3525 0.685 0.3525 0.82 0.205 0.82  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.04 0.36 0.155 0.36 0.155 0.52 0.35 0.52 0.35 0.485 0.415 0.485 0.415 0.62 0.35 0.62 0.35 0.585 0.14 0.585 0.14 1.12 0.04 1.12  ;
        POLYGON 0.48 0.36 0.545 0.36 0.545 0.745 0.95 0.745 0.95 0.71 1.015 0.71 1.015 0.845 0.95 0.845 0.95 0.81 0.545 0.81 0.545 0.98 0.48 0.98  ;
        POLYGON 1.28 0.81 1.315 0.81 1.315 0.595 0.86 0.595 0.86 0.53 1.38 0.53 1.38 0.81 1.415 0.81 1.415 0.875 1.28 0.875  ;
        POLYGON 0.655 0.875 0.72 0.875 0.72 1.005 1.48 1.005 1.48 0.43 1.365 0.43 1.365 0.465 1.3 0.465 1.3 0.33 1.365 0.33 1.365 0.365 1.545 0.365 1.545 0.935 2.35 0.935 2.35 1.145 2.285 1.145 2.285 1 1.58 1 1.58 1.21 1.515 1.21 1.515 1.07 0.72 1.07 0.72 1.15 0.655 1.15  ;
        POLYGON 1.61 0.655 2.23 0.655 2.23 0.4 2.16 0.4 2.16 0.335 2.295 0.335 2.295 0.665 2.48 0.665 2.48 0.835 2.515 0.835 2.515 1.11 2.45 1.11 2.45 0.97 2.415 0.97 2.415 0.73 2.26 0.73 2.26 0.72 1.61 0.72  ;
        POLYGON 2.36 0.495 2.885 0.495 2.885 0.56 2.36 0.56  ;
        POLYGON 3.08 0.495 3.215 0.495 3.215 0.535 3.845 0.535 3.845 0.88 3.915 0.88 3.915 0.945 3.78 0.945 3.78 0.6 3.155 0.6 3.155 0.56 3.08 0.56  ;
        POLYGON 2.735 0.935 2.955 0.935 2.955 0.97 3.585 0.97 3.585 1.04 4 1.04 4 0.93 4.325 0.93 4.325 1.02 4.555 1.02 4.555 0.945 4.52 0.945 4.52 0.88 4.555 0.88 4.555 0.685 4.11 0.685 4.11 0.55 4.175 0.55 4.175 0.62 4.62 0.62 4.62 0.88 4.655 0.88 4.655 0.945 4.62 0.945 4.62 1.085 4.26 1.085 4.26 0.995 4.065 0.995 4.065 1.105 3.52 1.105 3.52 1.035 2.855 1.035 2.855 1 2.67 1 2.67 0.625 2.95 0.625 2.95 0.335 3.165 0.335 3.165 0.4 3.015 0.4 3.015 0.69 2.735 0.69  ;
        POLYGON 4.415 1.15 4.72 1.15 4.72 0.295 4.41 0.295 4.41 0.33 4.345 0.33 4.345 0.295 4.15 0.295 4.15 0.23 4.345 0.23 4.345 0.195 4.41 0.195 4.41 0.23 4.785 0.23 4.785 1.215 4.415 1.215  ;
        POLYGON 4.85 0.32 4.915 0.32 4.915 0.5 5.465 0.5 5.4925 0.5 5.4925 0.465 5.5575 0.465 5.5575 0.6 5.4925 0.6 5.4925 0.565 5.465 0.565 5.1 0.565 5.1 0.76 5.035 0.76 5.035 0.565 4.85 0.565  ;
  END
END DFFRS_X2

MACRO DFFR_X1
  CLASS core ;
  FOREIGN DFFR_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.99 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.4825 0.5625 3.49 0.5625 3.49 0.4175 3.555 0.4175 3.555 1.115 3.49 1.115 3.49 0.6975 3.4825 0.6975  ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.435 0.4225 2.3425 0.4225 2.3425 0.15 2.86 0.15 2.86 0.4975 3.13 0.4975 3.13 0.5625 2.795 0.5625 2.795 0.215 2.4075 0.215 2.4075 0.4875 1.435 0.4875  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 0.8225 0.295 0.8225 0.295 1.315 0.555 1.315 0.555 1.0525 0.69 1.0525 0.69 1.315 1.38 1.315 1.38 1.0575 1.445 1.0575 1.445 1.315 2.15 1.315 2.15 0.9425 2.215 0.9425 2.215 1.315 2.92 1.315 2.92 1.0825 2.985 1.0825 2.985 1.315 3.315 1.315 3.315 1.0825 3.38 1.0825 3.38 1.315 3.675 1.315 3.675 1.04 3.74 1.04 3.74 1.315 3.99 1.315 3.99 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.8625 0.7025 3.865 0.7025 3.865 0.4175 3.93 0.4175 3.93 1.115 3.865 1.115 3.865 0.8375 3.8625 0.8375  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.095 0.2575 2.165 0.2575 2.165 0.085 1.65 0.085 1.65 0.3475 1.515 0.3475 1.515 0.2825 1.585 0.2825 1.585 0.085 0.69 0.085 0.69 0.2825 0.555 0.2825 0.555 0.2175 0.625 0.2175 0.625 0.085 0.3 0.085 0.3 0.3275 0.235 0.3275 0.235 0.085 0 0.085 0 -0.085 3.99 -0.085 3.99 0.085 3.74 0.085 3.74 0.5375 3.675 0.5375 3.675 0.085 3.025 0.085 3.025 0.4175 2.96 0.4175 2.96 0.085 2.23 0.085 2.23 0.3225 2.095 0.3225  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.5625 0.6975 0.5625 0.6975 0.6975 0.6325 0.6975  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.195 0.4225 0.3175 0.4225 0.3175 0.5575 0.195 0.5575  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.6625 0.05 0.6625 0.05 0.2975 0.115 0.2975 0.115 0.6225 0.37 0.6225 0.37 0.7575 0.305 0.7575 0.305 0.6875 0.11 0.6875 0.11 1.0425 0.045 1.0425  ;
        POLYGON 0.425 0.2975 0.49 0.2975 0.49 0.3975 0.5 0.3975 0.5 0.7775 0.86 0.7775 0.86 0.7075 0.925 0.7075 0.925 0.8425 0.5 0.8425 0.5 0.9575 0.435 0.9575 0.435 0.4325 0.425 0.4325  ;
        POLYGON 0.82 0.1675 1.215 0.1675 1.215 0.7475 1.15 0.7475 1.15 0.2325 0.885 0.2325 0.885 0.5475 0.82 0.5475  ;
        POLYGON 1.28 0.5525 1.93 0.5525 1.93 0.6175 1.28 0.6175  ;
        POLYGON 1.805 0.2225 2.01 0.2225 2.01 0.3575 1.805 0.3575  ;
        POLYGON 1.9 0.9425 2.01 0.9425 2.01 1.2175 1.945 1.2175 1.945 1.0775 1.9 1.0775  ;
        POLYGON 0.93 0.9075 1.02 0.9075 1.02 0.3625 0.95 0.3625 0.95 0.2975 1.085 0.2975 1.085 0.8125 2.125 0.8125 2.125 0.8775 1.825 0.8775 1.825 1.0875 1.76 1.0875 1.76 0.8775 1.085 0.8775 1.085 0.9725 0.995 0.9725 0.995 1.0475 1.065 1.0475 1.065 1.1125 0.93 1.1125  ;
        POLYGON 1.645 0.6825 2.47 0.6825 2.47 0.8175 2.405 0.8175 2.405 0.7475 1.645 0.7475  ;
        POLYGON 2.4725 0.4475 2.5375 0.4475 2.5375 0.5175 2.6 0.5175 2.6 0.7575 2.67 0.7575 2.67 0.8225 2.535 0.8225 2.535 0.5825 2.4725 0.5825  ;
        POLYGON 2.525 0.8875 2.735 0.8875 2.735 0.6925 2.665 0.6925 2.665 0.345 2.51 0.345 2.51 0.28 2.73 0.28 2.73 0.6275 3.205 0.6275 3.205 0.5575 3.27 0.5575 3.27 0.6925 2.8 0.6925 2.8 0.9525 2.59 0.9525 2.59 1.1625 2.525 1.1625  ;
        POLYGON 2.865 0.7575 2.93 0.7575 2.93 0.8275 3.335 0.8275 3.335 0.1975 3.4 0.1975 3.4 0.73 3.425 0.73 3.425 0.8925 3.175 0.8925 3.175 1.1625 3.11 1.1625 3.11 0.8925 2.865 0.8925  ;
  END
END DFFR_X1

MACRO DFFR_X2
  CLASS core ;
  FOREIGN DFFR_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.99 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.4825 0.7025 3.4875 0.7025 3.4875 0.3375 3.5525 0.3375 3.5525 1.1125 3.4875 1.1125 3.4875 0.8375 3.4825 0.8375  ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.4375 0.4225 2.3425 0.4225 2.3425 0.15 2.8625 0.15 2.8625 0.4975 3.1325 0.4975 3.1325 0.5625 2.7975 0.5625 2.7975 0.215 2.4075 0.215 2.4075 0.4875 1.4375 0.4875  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2325 1.315 0.2325 0.8225 0.2975 0.8225 0.2975 1.315 0.5575 1.315 0.5575 1.0525 0.6925 1.0525 0.6925 1.315 1.3825 1.315 1.3825 1.0575 1.4475 1.0575 1.4475 1.315 2.1525 1.315 2.1525 0.9425 2.2175 0.9425 2.2175 1.315 2.9225 1.315 2.9225 1.0825 2.9875 1.0825 2.9875 1.315 3.3175 1.315 3.3175 1.0825 3.3825 1.0825 3.3825 1.315 3.6725 1.315 3.6725 0.8925 3.7375 0.8925 3.7375 1.315 3.99 1.315 3.99 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.8625 0.3375 3.9275 0.3375 3.9275 1.1125 3.8625 1.1125  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.0925 0.2575 2.1625 0.2575 2.1625 0.085 1.6525 0.085 1.6525 0.3475 1.5175 0.3475 1.5175 0.2825 1.5875 0.2825 1.5875 0.085 0.6925 0.085 0.6925 0.2825 0.5575 0.2825 0.5575 0.2175 0.6275 0.2175 0.6275 0.085 0.3025 0.085 0.3025 0.3275 0.2375 0.3275 0.2375 0.085 0 0.085 0 -0.085 3.99 -0.085 3.99 0.085 3.7375 0.085 3.7375 0.3675 3.6725 0.3675 3.6725 0.085 3.0225 0.085 3.0225 0.4175 2.9575 0.4175 2.9575 0.085 2.2275 0.085 2.2275 0.3225 2.0925 0.3225  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.5625 0.6975 0.5625 0.6975 0.6975 0.6325 0.6975  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1975 0.4225 0.3175 0.4225 0.3175 0.5575 0.1975 0.5575  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.0475 0.6625 0.0525 0.6625 0.0525 0.2975 0.1175 0.2975 0.1175 0.6225 0.3725 0.6225 0.3725 0.7575 0.3075 0.7575 0.3075 0.6875 0.1125 0.6875 0.1125 1.0425 0.0475 1.0425  ;
        POLYGON 0.4275 0.2975 0.4925 0.2975 0.4925 0.3975 0.5025 0.3975 0.5025 0.7775 0.8625 0.7775 0.8625 0.7075 0.9275 0.7075 0.9275 0.8425 0.5025 0.8425 0.5025 0.9575 0.4375 0.9575 0.4375 0.4325 0.4275 0.4325  ;
        POLYGON 0.8225 0.1675 1.2175 0.1675 1.2175 0.7475 1.1525 0.7475 1.1525 0.2325 0.8875 0.2325 0.8875 0.5475 0.8225 0.5475  ;
        POLYGON 1.2825 0.5525 1.9275 0.5525 1.9275 0.6175 1.2825 0.6175  ;
        POLYGON 1.8025 0.2225 2.0075 0.2225 2.0075 0.3575 1.8025 0.3575  ;
        POLYGON 1.9025 0.9425 1.9675 0.9425 1.9675 1.0825 2.0125 1.0825 2.0125 1.2175 1.9025 1.2175  ;
        POLYGON 0.9325 0.9075 1.0225 0.9075 1.0225 0.3625 0.9525 0.3625 0.9525 0.2975 1.0875 0.2975 1.0875 0.8125 2.1275 0.8125 2.1275 0.8775 1.8275 0.8775 1.8275 1.0875 1.7625 1.0875 1.7625 0.8775 1.0875 0.8775 1.0875 0.9725 0.9975 0.9725 0.9975 1.0475 1.0675 1.0475 1.0675 1.1125 0.9325 1.1125  ;
        POLYGON 1.6425 0.6825 2.4725 0.6825 2.4725 0.8175 2.4075 0.8175 2.4075 0.7475 1.6425 0.7475  ;
        POLYGON 2.4725 0.4475 2.5375 0.4475 2.5375 0.5175 2.6025 0.5175 2.6025 0.7575 2.6725 0.7575 2.6725 0.8225 2.5375 0.8225 2.5375 0.5825 2.4725 0.5825  ;
        POLYGON 2.5275 0.8875 2.7375 0.8875 2.7375 0.6925 2.6675 0.6925 2.6675 0.345 2.5075 0.345 2.5075 0.28 2.7325 0.28 2.7325 0.6275 3.2475 0.6275 3.2475 0.7625 3.1825 0.7625 3.1825 0.6925 2.8025 0.6925 2.8025 0.9525 2.5925 0.9525 2.5925 1.1625 2.5275 1.1625  ;
        POLYGON 2.8675 0.765 2.9325 0.765 2.9325 0.835 3.3325 0.835 3.3325 0.1975 3.3975 0.1975 3.3975 0.9 3.1775 0.9 3.1775 1.1625 3.1125 1.1625 3.1125 0.9 2.8675 0.9  ;
  END
END DFFR_X2

MACRO DFFS_X1
  CLASS core ;
  FOREIGN DFFS_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 4.18 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.8275 0.7375 3.98 0.7375 3.98 0.4175 4.045 0.4175 4.045 1.1575 3.98 1.1575 3.98 0.8025 3.8275 0.8025  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.475 0.5975 2.455 0.5975 2.455 0.6625 1.475 0.6625  ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.26 1.315 0.26 1.0075 0.325 1.0075 0.325 1.315 0.62 1.315 0.62 1.0325 0.685 1.0325 0.685 1.315 1.43 1.315 1.43 1.1725 1.495 1.1725 1.495 1.315 2.215 1.315 2.215 1.2075 2.35 1.2075 2.35 1.315 2.97 1.315 2.97 1.1675 3.105 1.1675 3.105 1.315 3.79 1.315 3.79 1.0825 3.855 1.0825 3.855 1.315 4.18 1.315 4.18 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.4475 0.7375 3.585 0.7375 3.585 0.4175 3.67 0.4175 3.67 0.5525 3.65 0.5525 3.65 0.8875 3.585 0.8875 3.585 0.8025 3.4475 0.8025  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 4.18 -0.085 4.18 0.085 3.855 0.085 3.855 0.5375 3.79 0.5375 3.79 0.085 3.355 0.085 3.355 0.4475 3.29 0.4475 3.29 0.085 2.36 0.085 2.36 0.11 2.225 0.11 2.225 0.085 1.425 0.085 1.425 0.2575 1.36 0.2575 1.36 0.085 0.295 0.085 0.295 0.2575 0.23 0.2575 0.23 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.7025 0.725 0.7025 0.725 0.8375 0.6325 0.8375  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.205 0.8075 0.27 0.8075 0.27 0.8775 0.3525 0.8775 0.3525 0.9425 0.205 0.9425  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 1.27 0.4525 1.76 0.4525 1.76 0.28 1.825 0.28 1.825 0.5175 1.27 0.5175  ;
        POLYGON 1.295 0.8875 1.755 0.8875 1.755 1.0125 1.825 1.0125 1.825 1.0775 1.69 1.0775 1.69 0.9525 1.295 0.9525  ;
        POLYGON 0.935 1.1475 1.3 1.1475 1.3 1.0425 1.625 1.0425 1.625 1.1425 2.085 1.1425 2.085 1.0775 2.1675 1.0775 2.1675 1.0275 2.625 1.0275 2.625 1.0925 2.2325 1.0925 2.2325 1.1425 2.15 1.1425 2.15 1.2075 1.56 1.2075 1.56 1.1075 1.365 1.1075 1.365 1.2125 0.87 1.2125 0.87 0.9675 0.5325 0.9675 0.5325 1.1775 0.465 1.1775 0.465 0.9225 0.485 0.9225 0.485 0.4175 0.55 0.4175 0.55 0.9025 0.88 0.9025 0.88 0.8875 0.975 0.8875 0.975 0.5775 1.04 0.5775 1.04 0.9525 0.935 0.9525  ;
        POLYGON 2.02 0.175 2.665 0.175 2.665 0.24 2.02 0.24  ;
        POLYGON 1 1.0175 1.105 1.0175 1.105 0.5125 0.965 0.5125 0.965 0.28 1.03 0.28 1.03 0.4475 1.17 0.4475 1.17 0.7275 2.94 0.7275 2.94 0.7925 1.17 0.7925 1.17 1.0775 1.135 1.0775 1.135 1.0825 1 1.0825  ;
        POLYGON 2.0375 0.8775 2.94 0.8775 2.94 0.9425 2.1025 0.9425 2.1025 1.0125 2.0375 1.0125  ;
        POLYGON 0.045 0.2275 0.11 0.2275 0.11 0.5775 0.355 0.5775 0.355 0.2875 0.835 0.2875 0.835 0.15 1.26 0.15 1.26 0.3225 1.63 0.3225 1.63 0.15 1.955 0.15 1.955 0.305 2.73 0.305 2.73 0.2225 3.2 0.2225 3.2 0.5125 3.4 0.5125 3.4 0.6475 3.335 0.6475 3.335 0.5775 3.135 0.5775 3.135 0.2875 2.795 0.2875 2.795 0.365 2.755 0.365 2.755 0.37 1.89 0.37 1.89 0.215 1.695 0.215 1.695 0.3875 1.195 0.3875 1.195 0.215 0.9 0.215 0.9 0.4525 0.765 0.4525 0.765 0.3525 0.42 0.3525 0.42 0.6425 0.14 0.6425 0.14 1.2275 0.075 1.2275 0.075 0.6325 0.045 0.6325  ;
        POLYGON 2.595 1.1575 2.6875 1.1575 2.6875 1.1425 2.84 1.1425 2.84 1.0175 2.87 1.0175 2.87 1.0075 3.005 1.0075 3.005 0.5325 2.125 0.5325 2.125 0.4675 2.845 0.4675 2.845 0.4075 2.98 0.4075 2.98 0.4675 3.07 0.4675 3.07 1.0075 3.38 1.0075 3.38 0.9525 3.85 0.9525 3.85 0.8825 3.915 0.8825 3.915 1.0175 3.515 1.0175 3.515 1.2125 3.415 1.2125 3.415 1.0725 2.905 1.0725 2.905 1.2075 2.73 1.2075 2.73 1.2225 2.595 1.2225  ;
  END
END DFFS_X1

MACRO DFFS_X2
  CLASS core ;
  FOREIGN DFFS_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.99 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.6375 0.4575 3.8725 0.4575 3.8725 0.3 3.9375 0.3 3.9375 1.2275 3.8725 1.2275 3.8725 0.5225 3.6375 0.5225  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.4875 0.625 1.5475 0.625 1.5475 0.5975 1.6825 0.5975 1.6825 0.625 2.4125 0.625 2.4125 0.69 1.4875 0.69  ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2725 1.315 0.2725 1.0075 0.3375 1.0075 0.3375 1.315 0.6325 1.315 0.6325 1.04 0.6975 1.04 0.6975 1.315 1.4425 1.315 1.4425 1.18 1.5075 1.18 1.5075 1.315 2.1725 1.315 2.1725 1.215 2.3075 1.215 2.3075 1.315 2.9275 1.315 2.9275 1.195 3.0625 1.195 3.0625 1.315 3.6825 1.315 3.6825 1.0075 3.7475 1.0075 3.7475 1.315 3.99 1.315 3.99 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.4525 0.425 3.4975 0.425 3.4975 0.285 3.5625 0.285 3.5625 0.56 3.4525 0.56  ;
        POLYGON 3.4525 0.7925 3.54 0.7925 3.54 0.8775 3.7725 0.8775 3.7725 0.9425 3.5625 0.9425 3.5625 1.2275 3.4975 1.2275 3.4975 0.9275 3.4525 0.9275  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.99 -0.085 3.99 0.085 3.7475 0.085 3.7475 0.33 3.6825 0.33 3.6825 0.085 3.2825 0.085 3.2825 0.3925 3.2175 0.3925 3.2175 0.085 2.3525 0.085 2.3525 0.17 2.2175 0.17 2.2175 0.085 1.4375 0.085 1.4375 0.2575 1.3725 0.2575 1.3725 0.085 0.3075 0.085 0.3075 0.2575 0.2425 0.2575 0.2425 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.7125 0.5275 0.7775 0.5275 0.7775 0.5975 0.9225 0.5975 0.9225 0.6625 0.7125 0.6625  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.8075 0.2825 0.8075 0.2825 0.8775 0.3525 0.8775 0.3525 0.9425 0.2175 0.9425  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 1.2825 0.4525 1.7725 0.4525 1.7725 0.28 1.8375 0.28 1.8375 0.5175 1.2825 0.5175  ;
        POLYGON 1.3075 0.895 1.7675 0.895 1.7675 1.02 1.8375 1.02 1.8375 1.085 1.7025 1.085 1.7025 0.96 1.3075 0.96  ;
        POLYGON 0.9475 1.1525 1.3125 1.1525 1.3125 1.05 1.6375 1.05 1.6375 1.15 2.0425 1.15 2.0425 1.085 2.115 1.085 2.115 1.055 2.5825 1.055 2.5825 1.12 2.17 1.12 2.17 1.15 2.1075 1.15 2.1075 1.215 1.5725 1.215 1.5725 1.115 1.3775 1.115 1.3775 1.2175 0.8825 1.2175 0.8825 0.9575 0.5425 0.9575 0.5425 1.1775 0.4775 1.1775 0.4775 0.91 0.4975 0.91 0.4975 0.4175 0.5625 0.4175 0.5625 0.8925 0.9875 0.8925 0.9875 0.5825 1.0525 0.5825 1.0525 0.9575 0.9475 0.9575  ;
        POLYGON 2.0325 0.235 2.4775 0.235 2.4775 0.1675 2.6125 0.1675 2.6125 0.3 2.0325 0.3  ;
        POLYGON 1.0125 1.0225 1.1175 1.0225 1.1175 0.5175 0.98 0.5175 0.98 0.4725 0.9775 0.4725 0.9775 0.28 1.0425 0.28 1.0425 0.4525 1.1825 0.4525 1.1825 0.755 2.9175 0.755 2.9175 0.82 1.1825 0.82 1.1825 1.0825 1.1475 1.0825 1.1475 1.0875 1.0125 1.0875  ;
        POLYGON 1.995 0.885 2.06 0.885 2.06 0.905 2.9575 0.905 2.9575 0.97 2.06 0.97 2.06 1.02 1.995 1.02  ;
        POLYGON 0.0575 0.2275 0.1225 0.2275 0.1225 0.5775 0.3675 0.5775 0.3675 0.2875 0.8475 0.2875 0.8475 0.15 1.1725 0.15 1.1725 0.3225 1.6425 0.3225 1.6425 0.15 1.9675 0.15 1.9675 0.365 2.6775 0.365 2.6775 0.1675 3.0725 0.1675 3.0725 0.4575 3.3625 0.4575 3.3625 0.5225 3.0075 0.5225 3.0075 0.2325 2.7425 0.2325 2.7425 0.425 2.7025 0.425 2.7025 0.43 1.9025 0.43 1.9025 0.215 1.7075 0.215 1.7075 0.3875 1.1075 0.3875 1.1075 0.215 0.9125 0.215 0.9125 0.4525 0.7775 0.4525 0.7775 0.3525 0.4325 0.3525 0.4325 0.6425 0.1525 0.6425 0.1525 1.2275 0.0875 1.2275 0.0875 0.6325 0.0575 0.6325  ;
        POLYGON 2.5525 1.185 2.7975 1.185 2.7975 1.065 3.3225 1.065 3.3225 0.69 2.9075 0.69 2.9075 0.67 2.8775 0.67 2.8775 0.56 2.1125 0.56 2.1125 0.495 2.8075 0.495 2.8075 0.3075 2.9425 0.3075 2.9425 0.615 2.955 0.615 2.955 0.625 3.8075 0.625 3.8075 0.76 3.7425 0.76 3.7425 0.69 3.3875 0.69 3.3875 0.975 3.4075 0.975 3.4075 1.25 3.3425 1.25 3.3425 1.13 2.8625 1.13 2.8625 1.25 2.5525 1.25  ;
  END
END DFFS_X2

MACRO DFF_X1
  CLASS core ;
  FOREIGN DFF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.42 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.85 0.3375 2.985 0.3375 2.985 0.4575 3.0125 0.4575 3.0125 0.5225 2.915 0.5225 2.915 1.0025 2.85 1.0025  ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 0.9025 0.295 0.9025 0.295 1.315 0.88 1.315 0.88 1.13 0.945 1.13 0.945 1.315 1.655 1.315 1.655 1.2075 1.72 1.2075 1.72 1.315 2.58 1.315 2.58 1.23 2.51 1.23 2.51 1.165 2.645 1.165 2.645 1.315 3.11 1.315 3.11 0.9275 3.175 0.9275 3.175 1.315 3.42 1.315 3.42 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.0675 0.5975 3.295 0.5975 3.295 0.3375 3.36 0.3375 3.36 1.0025 3.295 1.0025 3.295 0.6625 3.0675 0.6625  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.36 0.2225 2.43 0.2225 2.43 0.085 1.735 0.085 1.735 0.2875 1.6 0.2875 1.6 0.2225 1.67 0.2225 1.67 0.085 0.94 0.085 0.94 0.3225 0.875 0.3225 0.875 0.085 0.295 0.085 0.295 0.4075 0.23 0.4075 0.23 0.085 0 0.085 0 -0.085 3.42 -0.085 3.42 0.085 3.17 0.085 3.17 0.4575 3.105 0.4575 3.105 0.085 2.495 0.085 2.495 0.2875 2.36 0.2875  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.7875 0.5975 0.965 0.5975 0.965 0.5475 1.03 0.5475 1.03 0.6825 0.965 0.6825 0.965 0.6625 0.7875 0.6625  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.7025 0.3175 0.7025 0.3175 0.8375 0.2525 0.8375 0.2525 0.7675 0.175 0.7675  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.3775 0.11 0.3775 0.11 0.5725 0.275 0.5725 0.275 0.5025 0.34 0.5025 0.34 0.6375 0.11 0.6375 0.11 1.0725 0.045 1.0725  ;
        POLYGON 0.535 0.3775 0.6 0.3775 0.6 0.4175 1.365 0.4175 1.365 0.5525 1.3 0.5525 1.3 0.4825 0.6 0.4825 0.6 0.9325 0.535 0.9325  ;
        POLYGON 0.47 0.9975 0.665 0.9975 0.665 0.765 0.685 0.765 0.685 0.7475 1.525 0.7475 1.525 0.8125 0.73 0.8125 0.73 1.115 0.76 1.115 0.76 1.25 0.665 1.25 0.665 1.0625 0.405 1.0625 0.405 0.2475 0.69 0.2475 0.69 0.1875 0.755 0.1875 0.755 0.3225 0.69 0.3225 0.69 0.3125 0.47 0.3125  ;
        POLYGON 0.795 0.925 0.86 0.925 0.86 0.995 1.075 0.995 1.075 1.0775 1.8 1.0775 1.8 1.1425 1.325 1.1425 1.325 1.25 1.26 1.25 1.26 1.1425 1.01 1.1425 1.01 1.06 0.795 1.06  ;
        POLYGON 1.26 0.2025 1.325 0.2025 1.325 0.2875 1.495 0.2875 1.495 0.3625 1.82 0.3625 1.82 0.4275 1.43 0.4275 1.43 0.3525 1.2825 0.3525 1.2825 0.3375 1.26 0.3375  ;
        POLYGON 1.385 0.8775 1.59 0.8775 1.59 0.6825 1.15 0.6825 1.15 0.5475 1.215 0.5475 1.215 0.6175 1.655 0.6175 1.655 0.8775 2.085 0.8775 2.085 0.5625 2.15 0.5625 2.15 0.9725 2.085 0.9725 2.085 0.9425 1.45 0.9425 1.45 1.0125 1.385 1.0125  ;
        POLYGON 2.02 0.2025 2.085 0.2025 2.085 0.4325 2.54 0.4325 2.54 0.4975 2.02 0.4975  ;
        POLYGON 2.17 1.035 2.59 1.035 2.59 0.965 2.655 0.965 2.655 1.1 2.235 1.1 2.235 1.25 2.17 1.25  ;
        POLYGON 2.43 0.6225 2.605 0.6225 2.605 0.2725 2.67 0.2725 2.67 0.835 2.785 0.835 2.785 1.0675 2.98 1.0675 2.98 0.7975 3.165 0.7975 3.165 0.7275 3.23 0.7275 3.23 0.8625 3.045 0.8625 3.045 1.1325 2.8 1.1325 2.8 1.25 2.735 1.25 2.735 1.11 2.72 1.11 2.72 0.9 2.605 0.9 2.605 0.6875 2.43 0.6875  ;
  END
END DFF_X1

MACRO DFF_X2
  CLASS core ;
  FOREIGN DFF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.42 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.7225 0.2825 2.805 0.2825 2.805 0.7475 2.74 0.7475 2.74 0.4175 2.7225 0.4175  ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 0.9325 0.295 0.9325 0.295 1.315 0.8925 1.315 0.8925 1.13 0.9575 1.13 0.9575 1.315 1.7925 1.315 1.7925 1.205 1.8575 1.205 1.8575 1.315 2.5925 1.315 2.5925 1.2275 2.5225 1.2275 2.5225 1.1625 2.6575 1.1625 2.6575 1.315 3 1.315 3 0.6675 3.065 0.6675 3.065 1.315 3.42 1.315 3.42 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.0675 0.3175 3.115 0.3175 3.115 0.2675 3.25 0.2675 3.25 0.8875 3.185 0.8875 3.185 0.4025 3.0675 0.4025  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.36 0.2175 2.43 0.2175 2.43 0.085 1.735 0.085 1.735 0.2825 1.6 0.2825 1.6 0.2175 1.67 0.2175 1.67 0.085 0.94 0.085 0.94 0.3175 0.875 0.3175 0.875 0.085 0.295 0.085 0.295 0.4075 0.23 0.4075 0.23 0.085 0 0.085 0 -0.085 3.42 -0.085 3.42 0.085 2.99 0.085 2.99 0.3125 2.925 0.3125 2.925 0.085 2.495 0.085 2.495 0.2825 2.36 0.2825  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.7875 0.5975 0.9775 0.5975 0.9775 0.5775 1.0425 0.5775 1.0425 0.7125 0.9775 0.7125 0.9775 0.6625 0.7875 0.6625  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.7025 0.3175 0.7025 0.3175 0.8375 0.2525 0.8375  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.3775 0.11 0.3775 0.11 0.5725 0.275 0.5725 0.275 0.5025 0.34 0.5025 0.34 0.6375 0.11 0.6375 0.11 1.1025 0.045 1.1025  ;
        POLYGON 0.535 0.3775 0.6 0.3775 0.6 0.4475 1.365 0.4475 1.365 0.5825 1.3 0.5825 1.3 0.5125 0.6 0.5125 0.6 0.9625 0.535 0.9625  ;
        POLYGON 0.47 1.0275 0.6775 1.0275 0.6775 0.795 0.6975 0.795 0.6975 0.7775 1.525 0.7775 1.525 0.8425 0.7425 0.8425 0.7425 1.115 0.7725 1.115 0.7725 1.25 0.6775 1.25 0.6775 1.0925 0.405 1.0925 0.405 0.2475 0.69 0.2475 0.69 0.1825 0.755 0.1825 0.755 0.3175 0.69 0.3175 0.69 0.3125 0.47 0.3125  ;
        POLYGON 0.8075 0.925 0.8725 0.925 0.8725 0.995 1.33 0.995 1.33 1.1075 1.6775 1.1075 1.6775 1.075 1.8125 1.075 1.8125 1.14 1.735 1.14 1.735 1.1725 1.3375 1.1725 1.3375 1.25 1.2725 1.25 1.2725 1.14 1.265 1.14 1.265 1.06 0.8075 1.06  ;
        POLYGON 1.26 0.1975 1.325 0.1975 1.325 0.3175 1.485 0.3175 1.485 0.3575 1.82 0.3575 1.82 0.4225 1.425 0.4225 1.425 0.3825 1.2825 0.3825 1.2825 0.3675 1.26 0.3675  ;
        POLYGON 1.4375 0.9075 1.59 0.9075 1.59 0.7125 1.15 0.7125 1.15 0.5775 1.215 0.5775 1.215 0.6475 1.655 0.6475 1.655 0.905 2.0975 0.905 2.0975 0.56 2.1625 0.56 2.1625 0.97 1.61 0.97 1.61 1.0425 1.4375 1.0425  ;
        POLYGON 2.02 0.1975 2.085 0.1975 2.085 0.3475 2.51 0.3475 2.51 0.3775 2.52 0.3775 2.52 0.57 2.455 0.57 2.455 0.4125 2.02 0.4125  ;
        POLYGON 2.1825 1.0325 2.6175 1.0325 2.6175 0.9625 2.6825 0.9625 2.6825 1.0975 2.2475 1.0975 2.2475 1.2475 2.1825 1.2475  ;
        POLYGON 2.4425 0.635 2.585 0.635 2.585 0.17 2.65 0.17 2.65 0.6475 2.675 0.6475 2.675 0.8125 2.87 0.8125 2.87 0.5375 3.01 0.5375 3.01 0.4675 3.075 0.4675 3.075 0.6025 2.935 0.6025 2.935 0.8775 2.8125 0.8775 2.8125 1.2475 2.7475 1.2475 2.7475 0.8775 2.61 0.8775 2.61 0.7 2.4425 0.7  ;
  END
END DFF_X2

MACRO DLH_X1
  CLASS core ;
  FOREIGN DLH_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.09 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2475 1.315 0.2475 0.8675 0.3125 0.8675 0.3125 1.315 0.6225 1.315 0.6225 1.065 0.6875 1.065 0.6875 1.315 1.3775 1.315 1.3775 1.065 1.4425 1.065 1.4425 1.315 1.72 1.315 1.72 1.065 1.785 1.065 1.785 1.315 2.09 1.315 2.09 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.925 0.4175 1.99 0.4175 1.99 0.6675 2.0275 0.6675 2.0275 0.8975 1.99 0.8975 1.99 0.92 1.99 1.055 1.925 1.055 1.925 0.92 1.925 0.8975 1.925 0.8025 1.925 0.7375 1.925 0.6675  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.09 -0.085 2.09 0.085 1.8 0.085 1.8 0.23 1.8 0.5375 1.735 0.5375 1.735 0.23 1.735 0.085 1.4625 0.085 1.4625 0.195 1.3975 0.195 1.3975 0.085 0.7075 0.085 0.7075 0.195 0.6425 0.195 0.6425 0.085 0.3125 0.085 0.3125 0.2125 0.2475 0.2125 0.2475 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.5975 0.4575 0.7225 0.4575 0.7225 0.29 0.7875 0.29 0.7875 0.4575 0.7875 0.5225 0.7325 0.5225 0.7325 0.7725 0.7325 0.8475 0.5975 0.8475 0.5975 0.7725  ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1925 0.5975 0.2575 0.5975 0.2575 0.7375 0.3525 0.7375 0.3525 0.8025 0.1925 0.8025  ;
    END
  END G
  OBS
      LAYER metal1 ;
        POLYGON 0.0625 0.1825 0.1275 0.1825 0.1275 0.3075 0.3575 0.3075 0.3575 0.4425 0.1275 0.4425 0.1275 0.9975 0.0625 0.9975  ;
        POLYGON 0.4375 0.7225 0.4675 0.7225 0.4675 0.3175 0.4375 0.3175 0.4375 0.1825 0.5025 0.1825 0.5025 0.2625 0.5325 0.2625 0.5325 0.9125 0.8725 0.9125 0.8725 0.895 0.8725 0.83 1.1425 0.83 1.1425 0.895 0.9375 0.895 0.9375 0.9775 0.8725 0.9775 0.5325 0.9775 0.5325 0.9975 0.4375 0.9975  ;
        POLYGON 1.0025 0.96 1.2075 0.96 1.2075 0.3 1.0225 0.3 1.0225 0.165 1.0875 0.165 1.0875 0.235 1.2075 0.235 1.21 0.235 1.2725 0.235 1.2725 0.8125 1.5225 0.8125 1.5225 0.8775 1.2725 0.8775 1.2725 1.025 1.0675 1.025 1.0675 1.235 1.0025 1.235  ;
        POLYGON 1.495 0.955 1.6 0.955 1.6 0.7475 1.4 0.7475 1.4 0.6125 1.465 0.6125 1.465 0.6825 1.55 0.6825 1.55 0.4175 1.615 0.4175 1.615 0.6825 1.665 0.6825 1.665 0.955 1.665 1.02 1.6 1.02 1.6 1.195 1.535 1.195 1.535 1.02 1.495 1.02  ;
  END
END DLH_X1

MACRO DLH_X2
  CLASS core ;
  FOREIGN DLH_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.09 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2325 1.315 0.2325 1.0075 0.2975 1.0075 0.2975 1.315 0.61 1.315 0.61 1.2075 0.675 1.2075 0.675 1.315 1.365 1.315 1.365 1.0675 1.43 1.0675 1.43 1.315 1.77 1.315 1.77 0.8675 1.835 0.8675 1.835 1.315 2.09 1.315 2.09 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.7375 0.7375 1.96 0.7375 1.96 0.4175 2.025 0.4175 2.025 1.0875 1.96 1.0875 1.96 0.8025 1.7375 0.8025  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.09 -0.085 2.09 0.085 1.835 0.085 1.835 0.4475 1.77 0.4475 1.77 0.085 1.495 0.085 1.495 0.2725 1.43 0.2725 1.43 0.085 0.74 0.085 0.74 0.2725 0.675 0.2725 0.675 0.085 0.295 0.085 0.295 0.33 0.23 0.33 0.23 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.55 0.2975 0.615 0.2975 0.615 0.3675 0.7325 0.3675 0.7325 0.905 0.6675 0.905 0.6675 0.5225 0.5975 0.5225 0.5975 0.4325 0.55 0.4325  ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1775 0.7375 0.2425 0.7375 0.2425 0.8775 0.3525 0.8775 0.3525 0.9425 0.1775 0.9425  ;
    END
  END G
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.3 0.11 0.3 0.11 0.5825 0.37 0.5825 0.37 0.7175 0.305 0.7175 0.305 0.6475 0.1125 0.6475 0.1125 1.1375 0.0475 1.1375 0.0475 0.6025 0.045 0.6025  ;
        POLYGON 0.4225 0.8625 0.465 0.8625 0.465 0.5575 0.43 0.5575 0.43 0.53 0.42 0.53 0.42 0.195 0.485 0.195 0.485 0.495 0.53 0.495 0.53 0.97 1.03 0.97 1.03 0.7975 1.095 0.7975 1.095 1.035 0.4875 1.035 0.4875 1.1375 0.4225 1.1375  ;
        POLYGON 0.955 1.1 1.16 1.1 1.16 0.7025 1.055 0.7025 1.055 0.2425 1.12 0.2425 1.12 0.6375 1.41 0.6375 1.41 0.5675 1.475 0.5675 1.475 0.7025 1.225 0.7025 1.225 1.165 0.955 1.165  ;
        POLYGON 1.325 0.3675 1.39 0.3675 1.39 0.4375 1.585 0.4375 1.585 0.4175 1.65 0.4175 1.65 0.9975 1.585 0.9975 1.585 0.5025 1.325 0.5025  ;
  END
END DLH_X2

MACRO DLL_X1
  CLASS core ;
  FOREIGN DLL_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.9 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 1.03 0.295 1.03 0.295 1.315 0.59 1.315 0.59 0.9425 0.655 0.9425 0.655 1.315 1.395 1.315 1.395 1.1825 1.325 1.1825 1.325 1.1175 1.46 1.1175 1.46 1.315 1.565 1.315 1.565 0.9125 1.63 0.9125 1.63 1.315 1.9 1.315 1.9 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.5825 0.5625 1.755 0.5625 1.755 0.3675 1.82 0.3675 1.82 1.0325 1.755 1.0325 1.755 0.6975 1.5825 0.6975  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.9 -0.085 1.9 0.085 1.63 0.085 1.63 0.4875 1.565 0.4875 1.565 0.085 1.41 0.085 1.41 0.3175 1.345 0.3175 1.345 0.085 0.655 0.085 0.655 0.3175 0.59 0.3175 0.59 0.085 0.31 0.085 0.31 0.2425 0.245 0.2425 0.245 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.4225 0.6975 0.4225 0.6975 0.5575 0.6325 0.5575  ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.205 0.7025 0.3175 0.7025 0.3175 0.8375 0.205 0.8375  ;
    END
  END GN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.43 0.06 0.43 0.06 0.2125 0.125 0.2125 0.125 0.4075 0.305 0.4075 0.305 0.3375 0.37 0.3375 0.37 0.4725 0.11 0.4725 0.11 1.25 0.045 1.25  ;
        POLYGON 0.435 0.2125 0.5 0.2125 0.5 0.6225 0.84 0.6225 0.84 0.5525 0.905 0.5525 0.905 0.6875 0.5 0.6875 0.5 1.1875 0.435 1.1875  ;
        POLYGON 0.965 0.7575 0.97 0.7575 0.97 0.1975 1.035 0.1975 1.035 0.6475 1.225 0.6475 1.225 0.7825 1.03 0.7825 1.03 1.1625 0.965 1.1625  ;
        POLYGON 1.41 0.9475 1.48 0.9475 1.48 1.0125 1.345 1.0125 1.345 0.8725 1.285 0.8725 1.285 0.8075 1.335 0.8075 1.335 0.3925 1.48 0.3925 1.48 0.4575 1.4 0.4575 1.4 0.8075 1.42 0.8075 1.42 0.8725 1.41 0.8725  ;
  END
END DLL_X1

MACRO DLL_X2
  CLASS core ;
  FOREIGN DLL_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.9 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 1.03 0.295 1.03 0.295 1.315 0.59 1.315 0.59 0.9425 0.655 0.9425 0.655 1.315 1.36 1.315 1.36 1.0825 1.425 1.0825 1.425 1.315 1.5875 1.315 1.5875 0.9375 1.6525 0.9375 1.6525 1.315 1.9 1.315 1.9 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.7725 0.3825 1.8375 0.3825 1.8375 1.1575 1.7725 1.1575  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.9 -0.085 1.9 0.085 1.6525 0.085 1.6525 0.4125 1.5875 0.4125 1.5875 0.085 1.425 0.085 1.425 0.3175 1.36 0.3175 1.36 0.085 0.655 0.085 0.655 0.3175 0.59 0.3175 0.59 0.085 0.31 0.085 0.31 0.2425 0.245 0.2425 0.245 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.4225 0.6975 0.4225 0.6975 0.4925 0.77 0.4925 0.77 0.5575 0.6325 0.5575  ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.17 0.7725 0.2525 0.7725 0.2525 0.7025 0.3175 0.7025 0.3175 0.8375 0.17 0.8375  ;
    END
  END GN
  OBS
      LAYER metal1 ;
        POLYGON 0.04 0.6125 0.045 0.6125 0.045 0.59 0.06 0.59 0.06 0.2125 0.125 0.2125 0.125 0.5025 0.355 0.5025 0.355 0.6375 0.105 0.6375 0.105 0.8625 0.11 0.8625 0.11 1.25 0.045 1.25 0.045 0.8875 0.04 0.8875  ;
        POLYGON 0.435 0.2125 0.5 0.2125 0.5 0.6225 0.92 0.6225 0.92 0.6875 0.5 0.6875 0.5 1.1875 0.435 1.1875  ;
        POLYGON 0.965 0.735 0.985 0.735 0.985 0.4225 0.965 0.4225 0.965 0.2875 1.05 0.2875 1.05 0.7175 1.3175 0.7175 1.3175 0.7825 1.03 0.7825 1.03 1.1625 0.965 1.1625  ;
        POLYGON 1.2075 0.9525 1.3825 0.9525 1.3825 0.6025 1.23 0.6025 1.23 0.5375 1.3825 0.5375 1.3825 0.3825 1.4475 0.3825 1.4475 1.0175 1.2075 1.0175  ;
  END
END DLL_X2

MACRO FA_X1
  CLASS core ;
  FOREIGN FA_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.42 BY 1.4 ;
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.285 0.24 3.385 0.24 3.385 1.085 3.285 1.085  ;
    END
  END S
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.555 0.5075 0.555 1.62 0.555 1.62 0.62 0.63 0.62 0.63 0.63 0.5075 0.63 0.5075 0.6975 0.4425 0.6975  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.745 1.315 3.095 1.315 3.095 1.01 3.16 1.01 3.16 1.315 3.42 1.315 3.42 1.485 0 1.485 0 1.315 0.285 1.315 0.285 0.975 0.35 0.975 0.35 1.315 1.035 1.315 1.035 1.075 1.17 1.075 1.17 1.14 1.1 1.14 1.1 1.315 1.415 1.315 1.415 1.075 1.48 1.075 1.48 1.315 2.68 1.315 2.68 1.11 2.815 1.11 2.815 1.175 2.745 1.175  ;
    END
  END VDD
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.4225 0.07 0.4225 0.07 0.15 0.17 0.15 0.17 1.05 0.07 1.05 0.07 0.5575 0.0625 0.5575  ;
    END
  END CO
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.42 -0.085 3.42 0.085 3.16 0.085 3.16 0.36 3.095 0.36 3.095 0.085 2.745 0.085 2.745 0.26 2.815 0.26 2.815 0.325 2.68 0.325 2.68 0.085 1.545 0.085 1.545 0.32 1.48 0.32 1.48 0.085 1.11 0.085 1.11 0.23 1.045 0.23 1.045 0.085 0.39 0.085 0.39 0.195 0.255 0.195 0.255 0.085 0 0.085  ;
    END
  END VSS
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.795 0.815 1.81 0.815 1.81 0.8 1.945 0.8 1.945 0.9325 1.945 0.9425 1.945 1.115 2.4 1.115 2.4 0.85 2.61 0.85 2.61 0.78 2.675 0.78 2.675 0.915 2.465 0.915 2.465 1.18 1.88 1.18 1.88 0.9425 1.7375 0.9425 1.7375 0.88 0.795 0.88  ;
    END
  END CI
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.365 0.425 1.75 0.425 1.75 0.4225 1.75 0.185 2.465 0.185 2.465 0.52 3.09 0.52 3.09 0.585 2.4 0.585 2.4 0.25 1.815 0.25 1.815 0.4225 1.8375 0.4225 1.8375 0.5575 1.75 0.5575 1.75 0.49 0.365 0.49  ;
    END
  END B
  OBS
      LAYER metal1 ;
        POLYGON 0.86 0.15 0.925 0.15 0.925 0.295 1.235 0.295 1.235 0.15 1.3 0.15 1.3 0.36 0.86 0.36  ;
        POLYGON 0.85 0.955 0.95 0.955 0.95 0.945 1.22 0.945 1.22 0.95 1.36 0.95 1.36 1.015 1.195 1.015 1.195 1.01 0.985 1.01 0.985 1.02 0.85 1.02  ;
        POLYGON 0.3 0.845 0.48 0.845 0.48 0.95 0.665 0.95 0.665 0.685 1.665 0.685 1.665 0.67 2.14 0.67 2.14 0.6 2.205 0.6 2.205 0.735 1.71 0.735 1.71 0.75 0.73 0.75 0.73 0.95 0.765 0.95 0.765 1.015 0.415 1.015 0.415 0.91 0.235 0.91 0.235 0.26 0.665 0.26 0.665 0.15 0.73 0.15 0.73 0.325 0.3 0.325  ;
        POLYGON 2.53 0.28 2.595 0.28 2.595 0.39 2.875 0.39 2.875 0.355 2.905 0.355 2.905 0.28 2.97 0.28 2.97 0.415 2.935 0.415 2.935 0.455 2.535 0.455 2.535 0.415 2.53 0.415  ;
        POLYGON 2.53 0.98 2.97 0.98 2.97 1.115 2.905 1.115 2.905 1.045 2.595 1.045 2.595 1.115 2.53 1.115  ;
        POLYGON 2.2 0.985 2.27 0.985 2.27 0.38 2.2 0.38 2.2 0.315 2.335 0.315 2.335 0.65 3.22 0.65 3.22 0.785 3.155 0.785 3.155 0.715 2.335 0.715 2.335 1.05 2.2 1.05  ;
  END
END FA_X1

MACRO FILLCELL_X1
  CLASS core ;
  FOREIGN FILLCELL_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.19 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.19 1.315 0.19 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.19 -0.085 0.19 0.085 0 0.085  ;
    END
  END VSS
END FILLCELL_X1

MACRO FILLCELL_X16
  CLASS core ;
  FOREIGN FILLCELL_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.04 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 3.04 1.315 3.04 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.04 -0.085 3.04 0.085 0 0.085  ;
    END
  END VSS
END FILLCELL_X16

MACRO FILLCELL_X2
  CLASS core ;
  FOREIGN FILLCELL_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0 0.085  ;
    END
  END VSS
END FILLCELL_X2

MACRO FILLCELL_X32
  CLASS core ;
  FOREIGN FILLCELL_X32 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 6.08 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 6.08 1.315 6.08 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 6.08 -0.085 6.08 0.085 0 0.085  ;
    END
  END VSS
END FILLCELL_X32

MACRO FILLCELL_X4
  CLASS core ;
  FOREIGN FILLCELL_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0 0.085  ;
    END
  END VSS
END FILLCELL_X4

MACRO FILLCELL_X8
  CLASS core ;
  FOREIGN FILLCELL_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 0 0.085  ;
    END
  END VSS
END FILLCELL_X8

MACRO HA_X1
  CLASS core ;
  FOREIGN HA_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.09 BY 1.4 ;
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.31 0.9125 1.3925 0.9125 1.3925 0.7025 1.7575 0.7025 1.7575 0.4925 1.5725 0.4925 1.5725 0.2425 1.6375 0.2425 1.6375 0.4275 1.8225 0.4275 1.8225 0.7675 1.4575 0.7675 1.4575 0.9775 1.31 0.9775  ;
    END
  END S
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.4225 0.5075 0.4225 0.5075 0.4675 0.7175 0.4675 0.7175 0.1875 1.1125 0.1875 1.1125 0.4425 1.5075 0.4425 1.5075 0.5075 1.0475 0.5075 1.0475 0.2525 0.7825 0.2525 0.7825 0.5325 0.5075 0.5325 0.5075 0.5575 0.4425 0.5575  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.0475 1.315 0.0475 0.915 0.1125 0.915 0.1125 1.315 0.4225 1.315 0.4225 0.915 0.4875 0.915 0.4875 1.315 1.795 1.315 1.795 0.9825 1.86 0.9825 1.86 1.315 2.09 1.315 2.09 1.485 0 1.485  ;
    END
  END VDD
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.98 0.95 1.9925 0.95 1.9925 0.6975 1.9475 0.6975 1.9475 0.2425 2.0275 0.2425 2.0275 0.6425 2.0575 0.6425 2.0575 0.95 2.0575 1.085 1.98 1.085  ;
    END
  END CO
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.09 -0.085 2.09 0.085 1.8225 0.085 1.8225 0.3625 1.7575 0.3625 1.7575 0.085 1.2425 0.085 1.2425 0.3625 1.1775 0.3625 1.1775 0.085 0.6525 0.085 0.6525 0.4025 0.5875 0.4025 0.5875 0.085 0.1125 0.085 0.1125 0.3575 0.0475 0.3575 0.0475 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1925 0.5525 0.2575 0.5525 0.2575 0.6225 0.7475 0.6225 0.7475 0.7575 0.6825 0.7575 0.6825 0.6875 0.1925 0.6875  ;
        POLYGON 1.2025 0.7025 1.2675 0.7025 1.2675 0.8375 1.2025 0.8375  ;
    END
  END B
  OBS
      LAYER metal1 ;
        POLYGON 1.16 0.9725 1.225 0.9725 1.225 1.0425 1.535 1.0425 1.535 0.9725 1.6 0.9725 1.6 1.1075 1.16 1.1075  ;
        POLYGON 0.9775 0.5725 1.6925 0.5725 1.6925 0.6375 0.9775 0.6375 0.9775 0.8825 0.9125 0.8825 0.9125 0.3825 0.8475 0.3825 0.8475 0.3175 0.9825 0.3175 0.9825 0.3825 0.9775 0.3825  ;
        POLYGON 0.1275 0.7525 0.29 0.7525 0.29 0.785 0.6175 0.785 0.6175 1.1725 1.5175 1.1725 1.53 1.1725 1.665 1.1725 1.665 0.8325 1.7975 0.8325 1.9275 0.8325 1.9275 0.8975 1.7975 0.8975 1.73 0.8975 1.73 1.2375 1.53 1.2375 1.5175 1.2375 0.5525 1.2375 0.5525 0.85 0.2975 0.85 0.2975 0.99 0.2325 0.99 0.2325 0.8175 0.07 0.8175 0.07 0.785 0.0625 0.785 0.0625 0.455 0.07 0.455 0.07 0.4225 0.3125 0.4225 0.3125 0.2925 0.5225 0.2925 0.5225 0.3575 0.3775 0.3575 0.3775 0.4875 0.1275 0.4875  ;
  END
END HA_X1

MACRO INV_X1
  CLASS core ;
  FOREIGN INV_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.7025 0.1275 0.7025 0.1275 0.8375 0.0625 0.8375  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 0.9025 0.11 0.9025 0.11 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0.11 0.085 0.11 0.3575 0.045 0.3575 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.4225 0.23 0.4225 0.23 0.2375 0.295 0.2375 0.295 0.9775 0.23 0.9775 0.23 0.5575 0.0625 0.5575  ;
    END
  END ZN
END INV_X1

MACRO INV_X16
  CLASS core ;
  FOREIGN INV_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.5925 0.1275 0.5925 0.1275 0.9775 0.0625 0.9775  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.0425 0.11 1.0425 0.11 1.315 0.42 1.315 0.42 1.0425 0.485 1.0425 0.485 1.315 0.8 1.315 0.8 1.0425 0.865 1.0425 0.865 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.865 0.085 0.865 0.4075 0.8 0.4075 0.8 0.085 0.485 0.085 0.485 0.4075 0.42 0.4075 0.42 0.085 0.11 0.085 0.11 0.4075 0.045 0.4075 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.2775 0.3 0.2775 0.3 0.5975 0.61 0.5975 0.61 0.2775 0.675 0.2775 0.675 0.9925 0.61 0.9925 0.61 0.6625 0.3 0.6625 0.3 0.9925 0.235 0.9925  ;
    END
  END ZN
END INV_X16

MACRO INV_X2
  CLASS core ;
  FOREIGN INV_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.5625 0.1275 0.5625 0.1275 0.6975 0.0625 0.6975  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 0.7625 0.11 0.7625 0.11 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0.11 0.085 0.11 0.2175 0.045 0.2175 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.2825 0.23 0.2825 0.23 0.1875 0.295 0.1875 0.295 0.9825 0.23 0.9825 0.23 0.4175 0.0625 0.4175  ;
    END
  END ZN
END INV_X2

MACRO INV_X32
  CLASS core ;
  FOREIGN INV_X32 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.4575 0.1625 0.4575 0.1625 0.5225 0.1275 0.5225 0.1275 0.8375 0.0625 0.8375  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.0675 0.11 1.0675 0.11 1.315 0.42 1.315 0.42 1.0675 0.485 1.0675 0.485 1.315 0.8 1.315 0.8 1.0675 0.865 1.0675 0.865 1.315 1.18 1.315 1.18 1.0675 1.245 1.0675 1.245 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.52 -0.085 1.52 0.085 1.245 0.085 1.245 0.3525 1.18 0.3525 1.18 0.085 0.865 0.085 0.865 0.3525 0.8 0.3525 0.8 0.085 0.485 0.085 0.485 0.3525 0.42 0.3525 0.42 0.085 0.11 0.085 0.11 0.3525 0.045 0.3525 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3 0.8775 0.61 0.8775 0.61 0.6675 0.675 0.6675 0.675 0.8775 0.99 0.8775 0.99 0.6675 1.055 0.6675 1.055 0.8775 1.37 0.8775 1.37 0.6675 1.435 0.6675 1.435 0.9425 0.235 0.9425 0.235 0.275 0.3 0.275 0.3 0.4175 0.61 0.4175 0.61 0.275 0.675 0.275 0.675 0.485 0.99 0.485 0.99 0.275 1.055 0.275 1.055 0.485 1.37 0.485 1.37 0.275 1.435 0.275 1.435 0.55 0.61 0.55 0.61 0.4825 0.3 0.4825  ;
    END
  END ZN
END INV_X32

MACRO INV_X4
  CLASS core ;
  FOREIGN INV_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.4225 0.1275 0.4225 0.1275 0.6025 0.0625 0.6025  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.0425 0.11 1.0425 0.11 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0.11 0.085 0.11 0.3325 0.045 0.3325 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.8425 0.23 0.8425 0.23 0.2025 0.295 0.2025 0.295 0.9925 0.23 0.9925 0.23 0.9775 0.0625 0.9775  ;
    END
  END ZN
END INV_X4

MACRO INV_X8
  CLASS core ;
  FOREIGN INV_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.4225 0.1275 0.4225 0.1275 0.7375 0.1625 0.7375 0.1625 0.8025 0.0625 0.8025  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 0.9925 0.11 0.9925 0.11 1.315 0.42 1.315 0.42 0.9925 0.485 0.9925 0.485 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.485 0.085 0.485 0.3575 0.42 0.3575 0.42 0.085 0.11 0.085 0.11 0.3575 0.045 0.3575 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.8775 0.23 0.8775 0.23 0.2275 0.295 0.2275 0.295 0.8775 0.3525 0.8775 0.3525 0.9425 0.2175 0.9425  ;
    END
  END ZN
END INV_X8

MACRO LOGIC0_X1
  CLASS core ;
  FOREIGN LOGIC0_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.2825 0.1575 0.2825 0.1575 0.4175 0.0625 0.4175  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.0925 1.315 0.0925 1.115 0.1575 1.115 0.1575 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0.1575 0.085 0.1575 0.2175 0.0925 0.2175 0.0925 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.1075 0.635 0.1725 0.635 0.1725 1.05 0.1075 1.05  ;
  END
END LOGIC0_X1

MACRO LOGIC1_X1
  CLASS core ;
  FOREIGN LOGIC1_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.38 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.8425 0.1575 0.8425 0.1575 1.1175 0.0625 1.1175  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.1375 1.315 0.1375 1.1825 0.2025 1.1825 0.2025 1.315 0.38 1.315 0.38 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.38 -0.085 0.38 0.085 0.2025 0.085 0.2025 0.145 0.1375 0.145 0.1375 0.085 0 0.085  ;
    END
  END VSS
  OBS
      LAYER metal1 ;
        POLYGON 0.1525 0.21 0.2575 0.21 0.2575 0.485 0.1525 0.485  ;
  END
END LOGIC1_X1

MACRO MUX2_X1
  CLASS core ;
  FOREIGN MUX2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.2025 0.15 1.2675 0.15 1.2675 1.25 1.2025 1.25  ;
    END
  END Z
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1975 0.4225 0.3175 0.4225 0.3175 0.5575 0.1975 0.5575  ;
    END
  END S
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.5775 0.35 0.6425 0.35 0.6425 0.825 0.9075 0.825 0.9075 0.755 1.0125 0.755 1.0125 0.2825 1.0775 0.2825 1.0775 0.82 0.9725 0.82 0.9725 0.89 0.5775 0.89  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2375 1.315 0.2375 1.0825 0.3025 1.0825 0.3025 1.315 1.0125 1.315 1.0125 1.17 1.0775 1.17 1.0775 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 1.0625 0.085 1.0625 0.1925 0.9975 0.1925 0.9975 0.085 0.3025 0.085 0.3025 0.1925 0.2375 0.1925 0.2375 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.7775 0.4225 0.8875 0.4225 0.8875 0.5575 0.8425 0.5575 0.8425 0.76 0.7775 0.76  ;
    END
  END B
  OBS
      LAYER metal1 ;
        POLYGON 0.0525 0.1625 0.1175 0.1625 0.1175 0.6225 0.3825 0.6225 0.3825 0.7575 0.3175 0.7575 0.3175 0.6875 0.1175 0.6875 0.1175 1.1125 0.0525 1.1125  ;
        POLYGON 0.3925 1.1175 0.5275 1.1175 0.5275 1.185 0.7925 1.185 0.7925 1.115 0.9275 1.115 0.9275 1.18 0.8575 1.18 0.8575 1.25 0.4625 1.25 0.4625 1.1825 0.3925 1.1825  ;
        POLYGON 0.5125 0.985 1.0725 0.985 1.0725 0.915 1.1375 0.915 1.1375 1.05 0.7275 1.05 0.7275 1.12 0.5925 1.12 0.5925 1.05 0.4575 1.05 0.4575 1.02 0.4475 1.02 0.4475 0.22 0.6175 0.22 0.6175 0.15 0.6825 0.15 0.6825 0.285 0.5125 0.285  ;
  END
END MUX2_X1

MACRO MUX2_X2
  CLASS core ;
  FOREIGN MUX2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.2025 0.15 1.2675 0.15 1.2675 1.25 1.2025 1.25  ;
    END
  END Z
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1975 0.4225 0.3175 0.4225 0.3175 0.5575 0.1975 0.5575  ;
    END
  END S
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.5775 0.35 0.6425 0.35 0.6425 0.825 0.9075 0.825 0.9075 0.755 1.0125 0.755 1.0125 0.2825 1.0775 0.2825 1.0775 0.82 0.9725 0.82 0.9725 0.89 0.5775 0.89  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2375 1.315 0.2375 1.0825 0.3025 1.0825 0.3025 1.315 1.0125 1.315 1.0125 1.17 1.0775 1.17 1.0775 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 1.0625 0.085 1.0625 0.1925 0.9975 0.1925 0.9975 0.085 0.3025 0.085 0.3025 0.1925 0.2375 0.1925 0.2375 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.7775 0.4225 0.8875 0.4225 0.8875 0.5575 0.8425 0.5575 0.8425 0.76 0.7775 0.76  ;
    END
  END B
  OBS
      LAYER metal1 ;
        POLYGON 0.0525 0.1625 0.1175 0.1625 0.1175 0.6225 0.3825 0.6225 0.3825 0.7575 0.3175 0.7575 0.3175 0.6875 0.1175 0.6875 0.1175 1.1125 0.0525 1.1125  ;
        POLYGON 0.3925 1.1175 0.5275 1.1175 0.5275 1.185 0.7925 1.185 0.7925 1.115 0.9275 1.115 0.9275 1.18 0.8575 1.18 0.8575 1.25 0.4625 1.25 0.4625 1.1825 0.3925 1.1825  ;
        POLYGON 0.5125 0.985 1.0725 0.985 1.0725 0.8875 1.1375 0.8875 1.1375 1.05 0.7275 1.05 0.7275 1.12 0.5925 1.12 0.5925 1.05 0.4575 1.05 0.4575 1.02 0.4475 1.02 0.4475 0.22 0.6175 0.22 0.6175 0.15 0.6825 0.15 0.6825 0.285 0.5125 0.285  ;
  END
END MUX2_X2

MACRO NAND2_X1
  CLASS core ;
  FOREIGN NAND2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 0.9025 0.11 0.9025 0.11 1.315 0.42 1.315 0.42 0.9025 0.485 0.9025 0.485 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.4225 0.34 0.4225 0.34 0.6375 0.2525 0.6375  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.11 0.085 0.11 0.4575 0.045 0.4575 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.7025 0.1275 0.7025 0.1275 0.8375 0.0625 0.8375  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.7025 0.42 0.7025 0.42 0.3775 0.485 0.3775 0.485 0.8375 0.3 0.8375 0.3 0.9775 0.235 0.9775  ;
    END
  END ZN
END NAND2_X1

MACRO NAND2_X2
  CLASS core ;
  FOREIGN NAND2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 0.9025 0.11 0.9025 0.11 1.315 0.42 1.315 0.42 0.9025 0.485 0.9025 0.485 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.4225 0.34 0.4225 0.34 0.6775 0.2525 0.6775  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.11 0.085 0.11 0.5075 0.045 0.5075 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.7025 0.1275 0.7025 0.1275 0.8375 0.0625 0.8375  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.7725 0.42 0.7725 0.42 0.2775 0.485 0.2775 0.485 0.8375 0.3175 0.8375 0.3175 1.1175 0.3 1.1175 0.3 1.1225 0.235 1.1225  ;
    END
  END ZN
END NAND2_X2

MACRO NAND2_X4
  CLASS core ;
  FOREIGN NAND2_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.0675 1.315 0.0675 0.9725 0.1325 0.9725 0.1325 1.315 0.4425 1.315 0.4425 0.9725 0.5075 0.9725 0.5075 1.315 0.8225 1.315 0.8225 0.9725 0.8875 0.9725 0.8875 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.5725 0.6425 0.6375 0.6425 0.6375 0.7125 0.8225 0.7125 0.8225 0.7025 0.8875 0.7025 0.8875 0.8375 0.8225 0.8375 0.8225 0.7775 0.5725 0.7775  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.8875 0.085 0.8875 0.4375 0.8225 0.4375 0.8225 0.085 0.1325 0.085 0.1325 0.4375 0.0675 0.4375 0.0675 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1975 0.2175 0.7575 0.2175 0.7575 0.6075 0.6925 0.6075 0.6925 0.4175 0.6325 0.4175 0.6325 0.2825 0.2625 0.2825 0.2625 0.6075 0.1975 0.6075  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2575 0.8525 0.2875 0.8525 0.2875 0.8425 0.4425 0.8425 0.4425 0.3475 0.5075 0.3475 0.5075 0.8425 0.6975 0.8425 0.6975 1.1925 0.6325 1.1925 0.6325 0.9075 0.3225 0.9075 0.3225 1.1925 0.2575 1.1925  ;
    END
  END ZN
END NAND2_X4

MACRO NAND3_X1
  CLASS core ;
  FOREIGN NAND3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.0425 0.11 1.0425 0.11 1.315 0.42 1.315 0.42 1.0425 0.485 1.0425 0.485 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.7025 0.1275 0.7025 0.1275 0.8375 0.0625 0.8375  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.5625 0.53 0.5625 0.53 0.6975 0.4425 0.6975  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.11 0.085 0.11 0.4575 0.045 0.4575 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.2825 0.34 0.2825 0.34 0.6775 0.2525 0.6775  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.9325 0.2525 0.9325 0.2525 0.8425 0.61 0.8425 0.61 0.4175 0.675 0.4175 0.675 1.1175 0.61 1.1175 0.61 0.9775 0.3 0.9775 0.3 1.1175 0.235 1.1175  ;
    END
  END ZN
END NAND3_X1

MACRO NAND3_X2
  CLASS core ;
  FOREIGN NAND3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 0.8925 0.11 0.8925 0.11 1.315 0.42 1.315 0.42 0.8925 0.485 0.8925 0.485 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.5625 0.1275 0.5625 0.1275 0.6975 0.0625 0.6975  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.2825 0.53 0.2825 0.53 0.6775 0.465 0.6775 0.465 0.4175 0.4425 0.4175  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.11 0.085 0.11 0.425 0.045 0.425 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.5625 0.34 0.5625 0.34 0.6975 0.2525 0.6975  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.7625 0.61 0.7625 0.61 0.2775 0.675 0.2775 0.675 1.1125 0.61 1.1125 0.61 0.8275 0.3175 0.8275 0.3175 1.1175 0.235 1.1175  ;
    END
  END ZN
END NAND3_X2

MACRO NAND3_X4
  CLASS core ;
  FOREIGN NAND3_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.0675 1.315 0.0675 0.9975 0.1325 0.9975 0.1325 1.315 0.4425 1.315 0.4425 0.9975 0.5075 0.9975 0.5075 1.315 0.8225 1.315 0.8225 0.9975 0.8875 0.9975 0.8875 1.315 1.2025 1.315 1.2025 0.9975 1.2675 0.9975 1.2675 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.5625 0.1975 0.5625 0.1975 0.1525 1.1375 0.1525 1.1375 0.6725 1.0725 0.6725 1.0725 0.2175 0.2625 0.2175 0.2625 0.6725 0.1275 0.6725 0.1275 0.6975 0.0625 0.6975  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.7625 0.5475 0.8275 0.5475 0.8275 0.7375 0.9225 0.7375 0.9225 0.8025 0.7625 0.8025  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 1.2675 0.085 1.2675 0.42 1.2025 0.42 1.2025 0.085 0.1325 0.085 0.1325 0.42 0.0675 0.42 0.0675 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4025 0.2825 0.9775 0.2825 0.9775 0.6725 0.9125 0.6725 0.9125 0.3475 0.5075 0.3475 0.5075 0.5575 0.4675 0.5575 0.4675 0.6725 0.4025 0.6725  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.8425 0.6325 0.8425 0.6325 0.4125 0.6975 0.4125 0.6975 0.8675 1.0125 0.8675 1.0125 0.7375 1.0775 0.7375 1.0775 1.0125 1.0125 1.0125 1.0125 0.9325 0.6975 0.9325 0.6975 0.9475 0.6325 0.9475 0.6325 0.9075 0.3175 0.9075 0.3175 1.1175 0.2525 1.1175  ;
    END
  END ZN
END NAND3_X4

MACRO NAND4_X1
  CLASS core ;
  FOREIGN NAND4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.0325 0.11 1.0325 0.11 1.315 0.42 1.315 0.42 1.0325 0.485 1.0325 0.485 1.315 0.8 1.315 0.8 1.0325 0.865 1.0325 0.865 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.4225 0.34 0.4225 0.34 0.6775 0.2525 0.6775  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.4225 0.72 0.4225 0.72 0.6775 0.6325 0.6775  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.11 0.085 0.11 0.5525 0.045 0.5525 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.7025 0.53 0.7025 0.53 0.8375 0.4425 0.8375  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.7025 0.1275 0.7025 0.1275 0.8375 0.0625 0.8375  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.9025 0.62 0.9025 0.62 0.8725 0.8 0.8725 0.8 0.2775 0.865 0.2775 0.865 0.5625 0.8875 0.5625 0.8875 0.6975 0.865 0.6975 0.865 0.9375 0.675 0.9375 0.675 1.1075 0.61 1.1075 0.61 0.9675 0.295 0.9675 0.295 1.1075 0.23 1.1075 0.23 1.0825 0.2175 1.0825  ;
    END
  END ZN
END NAND4_X1

MACRO NAND4_X2
  CLASS core ;
  FOREIGN NAND4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 0.8975 0.11 0.8975 0.11 1.315 0.42 1.315 0.42 0.8975 0.485 0.8975 0.485 1.315 0.8 1.315 0.8 0.8975 0.865 0.8975 0.865 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.5625 0.34 0.5625 0.34 0.6975 0.2525 0.6975  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.2825 0.72 0.2825 0.72 0.6775 0.655 0.6775 0.655 0.4175 0.6325 0.4175  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.11 0.085 0.11 0.335 0.045 0.335 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.2825 0.53 0.2825 0.53 0.6775 0.465 0.6775 0.465 0.4175 0.4425 0.4175  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.5625 0.1275 0.5625 0.1275 0.6975 0.0625 0.6975  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.7675 0.6225 0.7675 0.6225 0.7425 0.8 0.7425 0.8 0.2775 0.865 0.2775 0.865 0.8075 0.675 0.8075 0.675 1.1175 0.61 1.1175 0.61 0.8325 0.3175 0.8325 0.3175 1.1175 0.235 1.1175  ;
    END
  END ZN
END NAND4_X2

MACRO NAND4_X4
  CLASS core ;
  FOREIGN NAND4_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.71 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.0675 1.315 0.0675 1.0675 0.1325 1.0675 0.1325 1.315 0.4075 1.315 0.4075 1.2425 0.5425 1.2425 0.5425 1.315 0.7875 1.315 0.7875 1.2425 0.9225 1.2425 0.9225 1.315 1.1675 1.315 1.1675 1.2425 1.3025 1.2425 1.3025 1.315 1.5825 1.315 1.5825 1.0675 1.6475 1.0675 1.6475 1.315 1.71 1.315 1.71 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3625 0.52 0.4275 0.52 1.2875 0.52 1.3525 0.52 1.3525 0.8775 1.4925 0.8775 1.4925 0.9425 1.2875 0.9425 1.2875 0.585 0.4275 0.585 0.4275 0.7625 0.3625 0.7625  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.7425 0.7375 0.9225 0.7375 0.9225 0.8025 0.8075 0.8025 0.8075 0.8925 0.7425 0.8925 0.7425 0.8025  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.71 -0.085 1.71 0.085 1.6475 0.085 1.6475 0.335 1.5825 0.335 1.5825 0.085 0.1325 0.085 0.1325 0.195 0.0675 0.195 0.0675 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.8775 0.58 0.8775 0.58 0.9225 0.6175 0.9225 0.6525 0.9225 0.6525 0.9575 1.0975 0.9575 1.0975 0.8875 1.1625 0.8875 1.1625 1.0225 0.5175 1.0225 0.5175 0.9425 0.4075 0.9425  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2125 0.39 0.2775 0.39 1.0125 0.39 1.0125 0.2825 1.0775 0.2825 1.0775 0.39 1.4775 0.39 1.5425 0.39 1.5425 0.6775 1.4775 0.6775 1.4775 0.455 0.2775 0.455 0.2775 0.6775 0.2125 0.6775  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1475 0.81 0.3175 0.81 0.3175 1.0875 1.3925 1.0875 1.3925 1.0425 1.4575 1.0425 1.4575 1.1775 1.3925 1.1775 1.3925 1.155 1.0775 1.155 1.0775 1.2475 1.0125 1.2475 1.0125 1.1525 0.6975 1.1525 0.6975 1.2225 0.6325 1.2225 0.6325 1.1525 0.2525 1.1525 0.2525 0.875 0.0825 0.875 0.0825 0.26 0.1475 0.26 0.8225 0.26 0.8225 0.1575 0.8875 0.1575 0.8875 0.325 0.8225 0.325 0.1475 0.325  ;
    END
  END ZN
END NAND4_X4

MACRO NOR2_X1
  CLASS core ;
  FOREIGN NOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.09 0.11 1.09 0.11 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.7025 0.5075 0.7025 0.5075 0.8375 0.4425 0.8375  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.485 0.085 0.485 0.5375 0.42 0.5375 0.42 0.085 0.11 0.085 0.11 0.5375 0.045 0.5375 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.8425 0.1275 0.8425 0.1275 0.9775 0.0625 0.9775  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.4175 0.3 0.4175 0.3 0.9625 0.305 0.9625 0.305 0.9675 0.3125 0.9675 0.3125 0.9825 0.485 0.9825 0.485 1.1175 0.2525 1.1175 0.2525 1.0075 0.235 1.0075  ;
    END
  END ZN
END NOR2_X1

MACRO NOR2_X2
  CLASS core ;
  FOREIGN NOR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.57 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 0.8425 0.11 0.8425 0.11 1.315 0.57 1.315 0.57 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.4225 0.5075 0.4225 0.5075 0.5575 0.4425 0.5575  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.57 -0.085 0.57 0.085 0.485 0.085 0.485 0.3275 0.42 0.3275 0.42 0.085 0.11 0.085 0.11 0.3275 0.045 0.3275 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.4225 0.1275 0.4225 0.1275 0.5575 0.0625 0.5575  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.2975 0.3 0.2975 0.3 0.9825 0.42 0.9825 0.42 0.8425 0.485 0.8425 0.485 1.1175 0.2525 1.1175 0.2525 1.0275 0.235 1.0275  ;
    END
  END ZN
END NOR2_X2

MACRO NOR2_X4
  CLASS core ;
  FOREIGN NOR2_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.0525 1.315 0.0525 1.0225 0.1175 1.0225 0.1175 1.315 0.8075 1.315 0.8075 1.0225 0.8725 1.0225 0.8725 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.5625 0.5075 0.5625 0.5075 0.6975 0.4425 0.6975  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.5575 0.085 0.5575 0.3325 0.4925 0.3325 0.4925 0.085 0.1825 0.085 0.1825 0.3325 0.1175 0.3325 0.1175 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1825 0.7175 0.2475 0.7175 0.2475 1.1825 0.6325 1.1825 0.6325 0.8 0.6575 0.8 0.6575 0.7175 0.7275 0.7175 0.7275 0.8525 0.6975 0.8525 0.6975 1.2475 0.1825 1.2475  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3075 0.2025 0.3775 0.2025 0.3775 0.7625 0.4975 0.7625 0.4975 0.9825 0.5075 0.9825 0.5075 1.1175 0.4325 1.1175 0.4325 0.8275 0.3125 0.8275 0.3125 0.4775 0.3075 0.4775  ;
    END
  END ZN
END NOR2_X4

MACRO NOR3_X1
  CLASS core ;
  FOREIGN NOR3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 0.7625 0.11 0.7625 0.11 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.5625 0.1275 0.5625 0.1275 0.6975 0.0625 0.6975  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.5625 0.53 0.5625 0.53 0.6975 0.4425 0.6975  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.485 0.085 0.485 0.3675 0.42 0.3675 0.42 0.085 0.11 0.085 0.11 0.3675 0.045 0.3675 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.5925 0.34 0.5925 0.34 0.9775 0.2525 0.9775  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.2475 0.3 0.2475 0.3 0.4325 0.61 0.4325 0.61 0.2475 0.675 0.2475 0.675 0.5625 0.6975 0.5625 0.6975 0.6975 0.675 0.6975 0.675 0.9925 0.61 0.9925 0.61 0.4975 0.235 0.4975  ;
    END
  END ZN
END NOR3_X1

MACRO NOR3_X2
  CLASS core ;
  FOREIGN NOR3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 0.995 0.11 0.995 0.11 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.4225 0.1275 0.4225 0.1275 0.5875 0.0625 0.5875  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.8425 0.465 0.8425 0.465 0.5625 0.53 0.5625 0.53 0.9775 0.4425 0.9775  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.485 0.085 0.485 0.3575 0.42 0.3575 0.42 0.085 0.11 0.085 0.11 0.3575 0.045 0.3575 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.5625 0.34 0.5625 0.34 0.6975 0.2525 0.6975  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 1.1575 0.61 1.1575 0.61 0.4875 0.235 0.4875 0.235 0.3275 0.3 0.3275 0.3 0.4225 0.61 0.4225 0.61 0.3275 0.675 0.3275 0.675 0.5625 0.6975 0.5625 0.6975 0.6975 0.675 0.6975 0.675 1.2225 0.2175 1.2225  ;
    END
  END ZN
END NOR3_X2

MACRO NOR3_X4
  CLASS core ;
  FOREIGN NOR3_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.02 0.11 1.02 0.11 1.315 1.18 1.315 1.18 1.02 1.245 1.02 1.245 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.5875 0.24 0.5875 0.24 1.1825 1.0475 1.1825 1.0475 0.5225 0.9775 0.5225 0.9775 0.4575 1.1125 0.4575 1.1125 1.2475 0.175 1.2475  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.74 0.3175 0.9225 0.3175 0.9225 0.3825 0.805 0.3825 0.805 0.595 0.74 0.595  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 0.485 0.085 0.485 0.36 0.42 0.36 0.42 0.085 0.11 0.085 0.11 0.36 0.045 0.36 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.34 0.5875 0.405 0.5875 0.405 1.0525 0.7875 1.0525 0.7875 0.7375 0.87 0.7375 0.87 0.5875 0.935 0.5875 0.935 1.1175 0.34 1.1175  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.23 0.3 0.23 0.3 0.4575 0.61 0.4575 0.61 0.2175 0.675 0.2175 0.675 0.9875 0.61 0.9875 0.61 0.5225 0.235 0.5225  ;
    END
  END ZN
END NOR3_X4

MACRO NOR4_X1
  CLASS core ;
  FOREIGN NOR4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.085 1.315 0.085 0.9625 0.15 0.9625 0.15 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 1.1575 0.355 1.1575 0.355 0.7275 0.42 0.7275 0.42 1.2225 0.2175 1.2225  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.5975 1.1575 0.71 1.1575 0.71 0.7275 0.775 0.7275 0.775 1.2225 0.5975 1.2225  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.905 0.085 0.905 0.2975 0.84 0.2975 0.84 0.085 0.525 0.085 0.525 0.2975 0.46 0.2975 0.46 0.085 0.15 0.085 0.15 0.2975 0.085 0.2975 0.085 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.545 0.5975 0.7325 0.5975 0.7325 0.6625 0.61 0.6625 0.61 0.7325 0.545 0.7325  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.165 0.5975 0.3525 0.5975 0.3525 0.6625 0.23 0.6625 0.23 0.7325 0.165 0.7325  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.1775 0.3525 0.1775 0.3525 0.3625 0.65 0.3625 0.65 0.1775 0.715 0.1775 0.715 0.3925 0.905 0.3925 0.905 1.1275 0.84 1.1275 0.84 0.4575 0.66 0.4575 0.66 0.4275 0.275 0.4275 0.275 0.2425 0.2175 0.2425  ;
    END
  END ZN
END NOR4_X1

MACRO NOR4_X2
  CLASS core ;
  FOREIGN NOR4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.045 0.11 1.045 0.11 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.4225 0.34 0.4225 0.34 0.5575 0.2525 0.5575  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.7025 0.655 0.7025 0.655 0.4875 0.72 0.4875 0.72 0.8375 0.6325 0.8375  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.865 0.085 0.865 0.2275 0.8 0.2275 0.8 0.085 0.485 0.085 0.485 0.2275 0.42 0.2275 0.42 0.085 0.11 0.085 0.11 0.2275 0.045 0.2275 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.7025 0.465 0.7025 0.465 0.4875 0.53 0.4875 0.53 0.8375 0.4425 0.8375  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.4225 0.1275 0.4225 0.1275 0.5575 0.0625 0.5575  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.1775 0.295 0.1775 0.295 0.2925 0.61 0.2925 0.61 0.1975 0.675 0.1975 0.675 0.3225 0.865 0.3225 0.865 0.4225 0.8875 0.4225 0.8875 0.5575 0.865 0.5575 0.865 0.8875 0.8 0.8875 0.8 0.3875 0.62 0.3875 0.62 0.3575 0.2425 0.3575 0.2425 0.3325 0.23 0.3325 0.23 0.2425 0.2175 0.2425  ;
    END
  END ZN
END NOR4_X2

MACRO NOR4_X4
  CLASS core ;
  FOREIGN NOR4_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.71 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.05 1.315 0.05 1.2 0.185 1.2 0.185 1.315 1.6 1.315 1.6 1.06 1.665 1.06 1.665 1.315 1.71 1.315 1.71 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.5 0.81 1.25 0.81 1.25 0.535 1.395 0.535 1.395 0.6 1.315 0.6 1.315 0.81 1.315 0.875 0.435 0.875 0.435 0.81 0.435 0.6975 0.435 0.6 0.365 0.6 0.365 0.5625 0.365 0.535 0.5 0.535 0.5 0.5625 0.5075 0.5625 0.5075 0.6975 0.5 0.6975  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.77 0.36 0.7875 0.36 0.905 0.36 0.905 0.45 0.9225 0.45 0.9225 0.5225 0.7875 0.5225 0.7875 0.46 0.77 0.46  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.71 -0.085 1.71 0.085 1.665 0.085 1.665 0.2 1.6 0.2 1.6 0.085 1.325 0.085 1.325 0.165 1.19 0.165 1.19 0.085 0.945 0.085 0.945 0.165 0.81 0.165 0.81 0.085 0.565 0.085 0.565 0.165 0.43 0.165 0.43 0.085 0.185 0.085 0.185 0.165 0.05 0.165 0.05 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.665 0.68 1.085 0.68 1.085 0.49 1.15 0.49 1.15 0.745 1.085 0.745 0.665 0.745 0.6 0.745 0.6 0.5575 0.6 0.4225 0.6975 0.4225 0.6975 0.5575 0.665 0.5575  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.165 0.535 0.3 0.535 0.3 0.94 1.46 0.94 1.46 0.7025 1.495 0.7025 1.495 0.535 1.495 0.5 1.56 0.5 1.56 0.535 1.56 0.7025 1.665 0.7025 1.665 0.8375 1.525 0.8375 1.525 0.94 1.525 1.005 0.235 1.005 0.235 0.94 0.235 0.6 0.165 0.6  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.035 0.23 0.24 0.23 0.24 0.205 0.375 0.205 0.375 0.23 0.62 0.23 0.62 0.205 0.755 0.205 0.755 0.23 1 0.23 1 0.205 1.135 0.205 1.135 0.23 1.38 0.23 1.38 0.205 1.515 0.205 1.515 0.27 1.435 0.27 1.435 0.295 0.1 0.295 0.1 0.96 0.1 0.98 0.145 0.98 0.145 1.07 0.94 1.07 0.94 1.17 0.805 1.17 0.805 1.135 0.035 1.135 0.035 0.96  ;
    END
  END ZN
END NOR4_X4

MACRO OAI211_X1
  CLASS core ;
  FOREIGN OAI211_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.53 0.475 0.5975 0.475 0.5975 0.4575 0.7325 0.4575 0.7325 0.54 0.595 0.54 0.595 0.6475 0.53 0.6475  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.1475 0.11 1.1475 0.11 1.315 0.61 1.315 0.61 1.1475 0.675 1.1475 0.675 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.865 0.085 0.865 0.4275 0.8 0.4275 0.8 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.7025 0.72 0.7025 0.72 0.8375 0.6325 0.8375  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.235 0.3875 0.3 0.3875 0.3 1.0175 0.865 1.0175 0.865 1.2225 0.8 1.2225 0.8 1.0825 0.485 1.0825 0.485 1.2225 0.42 1.2225 0.42 1.0825 0.25 1.0825 0.25 1.06 0.235 1.06  ;
    END
  END ZN
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.5975 0.1625 0.5975 0.1625 0.6625 0.1275 0.6625 0.1275 0.8375 0.0625 0.8375  ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.365 0.6675 0.43 0.6675 0.43 0.7375 0.5425 0.7375 0.5425 0.8025 0.365 0.8025  ;
    END
  END C1
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.2575 0.485 0.2575 0.485 0.4275 0.42 0.4275 0.42 0.3225 0.11 0.3225 0.11 0.4275 0.045 0.4275  ;
  END
END OAI211_X1

MACRO OAI211_X2
  CLASS core ;
  FOREIGN OAI211_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.52 0.7825 0.59 0.7825 0.59 0.7375 0.655 0.7375 0.8875 0.7375 0.8875 0.8375 0.8225 0.8375 0.8225 0.8025 0.655 0.8025 0.655 0.8175 0.655 0.8475 0.52 0.8475  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.0675 0.11 1.0675 0.11 1.315 0.59 1.315 0.59 1.0425 0.725 1.0425 0.725 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.87 0.085 0.87 0.3925 0.805 0.3925 0.805 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.5975 0.4575 0.765 0.4575 0.765 0.545 0.835 0.545 0.835 0.61 0.7 0.61 0.7 0.5225 0.5975 0.5225  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2575 0.9125 0.88 0.9125 0.88 1.2275 0.815 1.2275 0.815 0.9775 0.52 0.9775 0.52 1.1275 0.385 1.1275 0.385 0.9775 0.2575 0.9775 0.1925 0.9775 0.1925 0.5625 0.1925 0.485 0.23 0.485 0.23 0.345 0.195 0.345 0.195 0.28 0.33 0.28 0.33 0.345 0.295 0.345 0.295 0.485 0.295 0.5625 0.2575 0.5625  ;
    END
  END ZN
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.7025 0.1275 0.7025 0.1275 0.8375 0.0625 0.8375  ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.35 0.5975 0.5425 0.5975 0.5425 0.6625 0.35 0.6625  ;
    END
  END C1
  OBS
      LAYER metal1 ;
        POLYGON 0.395 0.325 0.42 0.325 0.42 0.215 0.11 0.215 0.11 0.425 0.045 0.425 0.045 0.15 0.485 0.15 0.485 0.325 0.53 0.325 0.53 0.39 0.395 0.39  ;
  END
END OAI211_X2

MACRO OAI211_X4
  CLASS core ;
  FOREIGN OAI211_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.71 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.3925 0.7025 1.4125 0.7025 1.4125 0.5875 0.98 0.5875 0.98 0.6575 0.915 0.6575 0.915 0.5225 1.4775 0.5225 1.4775 0.8375 1.3925 0.8375  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.0675 0.11 1.0675 0.11 1.315 0.8 1.315 0.8 1.0675 0.865 1.0675 0.865 1.315 1.18 1.315 1.18 1.0675 1.245 1.0675 1.245 1.315 1.71 1.315 1.71 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.71 -0.085 1.71 0.085 1.28 0.085 1.28 0.3275 1.145 0.3275 1.145 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.065 0.6525 1.2675 0.6525 1.2675 0.8375 1.2025 0.8375 1.2025 0.7175 1.065 0.7175  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.425 0.9125 0.785 0.9125 0.785 0.5875 0.69 0.5875 0.69 0.585 0.6325 0.585 0.6325 0.555 0.295 0.555 0.295 0.455 0.2 0.455 0.2 0.39 0.335 0.39 0.335 0.4025 0.36 0.4025 0.36 0.49 0.575 0.49 0.575 0.39 0.71 0.39 0.71 0.5225 0.85 0.5225 0.85 0.9125 1.06 0.9125 1.06 0.9825 1.0775 0.9825 1.0775 1.1875 0.995 1.1875 0.995 0.9775 0.49 0.9775 0.49 1.1875 0.425 1.1875  ;
    END
  END ZN
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.5625 0.215 0.5625 0.215 0.6525 0.72 0.6525 0.72 0.7875 0.655 0.7875 0.655 0.7175 0.0625 0.7175  ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.7825 0.415 0.7825 0.415 0.8475 0.3175 0.8475 0.3175 1.1175 0.2525 1.1175  ;
    END
  END C1
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.215 0.11 0.215 0.11 0.26 0.425 0.26 0.425 0.15 0.49 0.15 0.49 0.1825 0.865 0.1825 0.865 0.3925 1.56 0.3925 1.56 0.1825 1.625 0.1825 1.625 0.4575 0.8 0.4575 0.8 0.2475 0.49 0.2475 0.49 0.425 0.425 0.425 0.425 0.325 0.11 0.325 0.11 0.49 0.045 0.49  ;
  END
END OAI211_X4

MACRO OAI21_X1
  CLASS core ;
  FOREIGN OAI21_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.7025 0.6975 0.7025 0.6975 0.84 0.6325 0.84  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.0625 1.315 0.0625 1.0425 0.1275 1.0425 0.1275 1.315 0.6275 1.315 0.6275 1.0425 0.6925 1.0425 0.6925 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3775 0.77 0.4425 0.77 0.4425 0.7025 0.51 0.7025 0.51 0.8375 0.4425 0.8375 0.4425 0.905 0.3775 0.905 0.3775 0.8375  ;
    END
  END B1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.6925 0.085 0.6925 0.4975 0.6275 0.4975 0.6275 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.795 0.1275 0.795 0.1275 0.9775 0.0625 0.9775  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2475 0.4175 0.3125 0.4175 0.3125 0.9825 0.5075 0.9825 0.5075 1.1175 0.4425 1.1175 0.4425 1.0475 0.2475 1.0475  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.0625 0.2875 0.5025 0.2875 0.5025 0.4975 0.4375 0.4975 0.4375 0.3525 0.1275 0.3525 0.1275 0.4975 0.0625 0.4975  ;
  END
END OAI21_X1

MACRO OAI21_X2
  CLASS core ;
  FOREIGN OAI21_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.8775 0.645 0.8775 0.645 0.9425 0.4075 0.9425  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.0675 0.11 1.0675 0.11 1.315 0.625 1.315 0.625 1.0675 0.69 1.0675 0.69 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.36 0.56 0.495 0.56 0.495 0.5975 0.5425 0.5975 0.5425 0.6625 0.4075 0.6625 0.4075 0.625 0.36 0.625  ;
    END
  END B1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.69 0.085 0.69 0.49 0.625 0.49 0.625 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1275 0.7975 0.1975 0.7975 0.1975 0.8625 0.0625 0.8625 0.0625 0.5975 0.1625 0.5975 0.1625 0.6625 0.1275 0.6625  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.295 0.6825 0.3275 0.6825 0.3275 1.0175 0.52 1.0175 0.52 1.2225 0.2175 1.2225 0.2175 1.1575 0.2625 1.1575 0.2625 0.74 0.23 0.74 0.23 0.5 0.195 0.5 0.195 0.295 0.33 0.295 0.33 0.5 0.295 0.5  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.405 0.39 0.42 0.39 0.42 0.23 0.11 0.23 0.11 0.49 0.045 0.49 0.045 0.165 0.485 0.165 0.485 0.39 0.54 0.39 0.54 0.455 0.405 0.455  ;
  END
END OAI21_X2

MACRO OAI21_X4
  CLASS core ;
  FOREIGN OAI21_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.875 0.6525 1.01 0.6525 1.01 0.7375 1.1125 0.7375 1.1125 0.8025 0.945 0.8025 0.945 0.7375 0.945 0.7175 0.875 0.7175  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.385 1.315 0.385 1.1025 0.52 1.1025 0.52 1.315 0.99 1.315 0.99 1.0675 1.055 1.0675 1.055 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.19 0.5975 0.6625 0.5975 0.665 0.5975 0.7275 0.5975 0.7275 0.6725 0.8 0.6725 0.8 0.7375 0.6625 0.7375 0.6625 0.6975 0.6625 0.6725 0.6625 0.6625 0.255 0.6625 0.255 0.7325 0.19 0.7325  ;
    END
  END B1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 1.095 0.085 1.095 0.4575 0.96 0.4575 0.96 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.305 0.7825 0.34 0.7825 0.4075 0.7825 0.4075 0.7375 0.5425 0.7375 0.5425 0.7825 0.5425 0.8025 0.475 0.8025 0.475 0.8475 0.34 0.8475 0.305 0.8475  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.11 0.8875 0.11 0.9125 0.865 0.9125 0.865 1.1875 0.8 1.1875 0.8 0.9775 0.1275 0.9775 0.1275 1.1175 0.11 1.1175 0.11 1.1625 0.045 1.1625 0.045 1.1175 0.045 0.8875 0.045 0.5025 0.045 0.4375 0.195 0.4375 0.195 0.3 0.195 0.2975 0.33 0.2975 0.33 0.3 0.33 0.4375 0.585 0.4375 0.585 0.2975 0.72 0.2975 0.72 0.5025 0.33 0.5025 0.32 0.5025 0.195 0.5025 0.11 0.5025  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.1675 0.11 0.1675 0.87 0.1675 0.87 0.5225 1.185 0.5225 1.185 0.2625 1.25 0.2625 1.25 0.5875 0.805 0.5875 0.805 0.2325 0.485 0.2325 0.485 0.3525 0.42 0.3525 0.42 0.2325 0.11 0.2325 0.11 0.3525 0.045 0.3525  ;
  END
END OAI21_X4

MACRO OAI221_X1
  CLASS core ;
  FOREIGN OAI221_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.5625 0.595 0.5625 0.595 0.6975 0.4425 0.6975  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.1725 0.11 1.1725 0.11 1.315 0.61 1.315 0.61 1.1725 0.675 1.1725 0.675 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.8425 0.34 0.8425 0.34 0.9775 0.2525 0.9775  ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.425 1.0425 0.805 1.0425 0.805 0.3275 0.87 0.3275 0.87 0.7025 0.8875 0.7025 0.8875 1.05 1.055 1.05 1.055 1.185 0.99 1.185 0.99 1.115 0.855 1.115 0.855 1.1075 0.49 1.1075 0.49 1.2475 0.425 1.2475  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.935 0.5225 1 0.5225 1 0.5625 1.0775 0.5625 1.0775 0.6975 1.0125 0.6975 1.0125 0.6575 0.935 0.6575  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.295 0.085 0.295 0.3675 0.23 0.3675 0.23 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.5625 0.1275 0.5625 0.1275 0.6975 0.0625 0.6975  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.8425 0.72 0.8425 0.72 0.9775 0.6325 0.9775  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.3275 0.11 0.3275 0.11 0.4325 0.42 0.4325 0.42 0.3275 0.485 0.3275 0.485 0.4625 0.48 0.4625 0.48 0.4975 0.045 0.4975  ;
        POLYGON 0.615 0.1975 1.055 0.1975 1.055 0.3675 0.99 0.3675 0.99 0.2625 0.68 0.2625 0.68 0.3675 0.615 0.3675  ;
  END
END OAI221_X1

MACRO OAI221_X2
  CLASS core ;
  FOREIGN OAI221_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.51 0.7425 0.6325 0.7425 0.6325 0.7025 0.6975 0.7025 0.6975 0.8375 0.51 0.8375  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.07 1.315 0.07 1.0075 0.135 1.0075 0.135 1.315 0.615 1.315 0.615 1.0425 0.75 1.0425 0.75 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.305 0.6875 0.375 0.6875 0.375 0.5975 0.5425 0.5975 0.5425 0.6625 0.44 0.6625 0.44 0.7525 0.305 0.7525  ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.91 0.9025 1.095 0.9025 1.095 1.1775 1.03 1.1775 1.03 0.9675 0.88 0.9675 0.88 0.9775 0.545 0.9775 0.545 1.1175 0.41 1.1175 0.41 0.9125 0.845 0.9125 0.845 0.345 0.81 0.345 0.81 0.28 0.945 0.28 0.945 0.345 0.91 0.345  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.0125 0.7025 1.0775 0.7025 1.0775 0.8375 1.0125 0.8375  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.32 0.085 0.32 0.3925 0.255 0.3925 0.255 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.5875 0.25 0.5875 0.25 0.6525 0.1275 0.6525 0.1275 0.8375 0.0625 0.8375  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.4225 0.6975 0.4225 0.6975 0.545 0.78 0.545 0.78 0.61 0.6325 0.61  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.07 0.245 0.135 0.245 0.135 0.4575 0.445 0.4575 0.445 0.245 0.51 0.245 0.51 0.5225 0.115 0.5225 0.115 0.52 0.07 0.52  ;
        POLYGON 0.61 0.1525 0.725 0.1525 0.725 0.15 1.095 0.15 1.095 0.425 1.03 0.425 1.03 0.215 0.745 0.215 0.745 0.3575 0.61 0.3575  ;
  END
END OAI221_X2

MACRO OAI221_X4
  CLASS core ;
  FOREIGN OAI221_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.28 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.0125 0.6525 1.2 0.6525 1.2 0.7175 1.0775 0.7175 1.0775 0.8375 1.0125 0.8375  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.405 1.315 0.405 1.1025 0.54 1.1025 0.54 1.315 1.145 1.315 1.145 1.1025 1.28 1.1025 1.28 1.315 2.055 1.315 2.055 1.1025 2.19 1.1025 2.19 1.315 2.28 1.315 2.28 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.785 0.7975 2.0275 0.7975 2.0275 0.9775 1.9625 0.9775 1.9625 0.8625 1.785 0.8625  ;
    END
  END B1
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.11 0.9725 1.81 0.9725 1.81 1.1775 1.675 1.1775 1.675 1.0375 0.11 1.0375 0.11 1.1625 0.045 1.1625 0.045 0.2775 0.13 0.2775 0.13 0.35 0.405 0.35 0.405 0.3125 0.54 0.3125 0.54 0.35 0.785 0.35 0.785 0.28 0.92 0.28 0.92 0.5225 0.805 0.5225 0.805 0.415 0.11 0.415  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.5875 0.815 0.5875 0.815 0.6525 0.6975 0.6525 0.6975 0.8375 0.6325 0.8375 0.6325 0.6525 0.175 0.6525  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.28 -0.085 2.28 0.085 2.03 0.085 2.03 0.425 1.965 0.425 1.965 0.085 1.65 0.085 1.65 0.425 1.585 0.425 1.585 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.445 0.6675 2.11 0.6675 2.11 0.7325 1.6475 0.7325 1.6475 0.8375 1.5825 0.8375 1.5825 0.7325 1.445 0.7325  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.7375 0.3925 0.7375 0.3925 0.7975 0.46 0.7975 0.46 0.8625 0.3525 0.8625 0.325 0.8625 0.325 0.8025 0.2175 0.8025  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.255 0.15 1.27 0.15 1.27 0.425 1.205 0.425 1.205 0.215 0.695 0.215 0.695 0.285 0.63 0.285 0.63 0.215 0.32 0.215 0.32 0.285 0.255 0.285  ;
        POLYGON 0.985 0.3125 1.12 0.3125 1.12 0.49 1.395 0.49 1.395 0.2775 1.46 0.2775 1.46 0.49 1.775 0.49 1.775 0.2775 1.84 0.2775 1.84 0.49 2.155 0.49 2.155 0.2775 2.22 0.2775 2.22 0.555 1.1 0.555 1.1 0.5525 0.985 0.5525  ;
  END
END OAI221_X4

MACRO OAI222_X1
  CLASS core ;
  FOREIGN OAI222_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2625 1.315 0.2625 1.1075 0.3275 1.1075 0.3275 1.315 1.3625 1.315 1.3625 1.025 1.4275 1.025 1.4275 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.7025 0.6975 0.7025 0.7525 0.7025 0.7525 0.8375 0.6975 0.8375 0.6325 0.8375  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.8225 0.7025 0.8875 0.7025 1.0025 0.7025 1.0025 0.8375 1.0025 0.9125 0.9375 0.9125 0.9375 0.8375 0.8875 0.8375 0.8225 0.8375  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.2025 0.5625 1.2675 0.5625 1.2675 0.6975 1.2025 0.6975  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6475 1.1075 0.7125 1.1075 0.7125 1.185 0.9875 1.185 0.9875 0.9775 1.0725 0.9775 1.0725 0.51 1.0475 0.51 1.0475 0.3225 1.0725 0.3225 1.1125 0.3225 1.1125 0.4575 1.1375 0.4575 1.1375 0.8425 1.2675 0.8425 1.2675 0.9775 1.1375 0.9775 1.1375 1.0425 1.0525 1.0425 1.0525 1.25 0.6475 1.25  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.7025 0.5075 0.7025 0.5625 0.7025 0.5625 0.8375 0.5075 0.8375 0.4425 0.8375  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4225 0.2625 0.4575 0.2625 0.4575 0.085 0 0.085 0 -0.085 1.52 -0.085 1.52 0.085 0.5225 0.085 0.5225 0.2625 0.5575 0.2625 0.5575 0.3275 0.5225 0.3275 0.4575 0.3275 0.4225 0.3275  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.7025 0.1275 0.7025 0.1275 0.8375 0.0625 0.8375  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.7025 0.3725 0.7025 0.3725 0.8375 0.2525 0.8375  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.2675 0.2475 0.3325 0.2475 0.3325 0.3925 0.6425 0.3925 0.6425 0.25 0.7075 0.25 0.7075 0.3925 0.7075 0.4275 0.7075 0.4575 0.2675 0.4575 0.2675 0.4275 0.2675 0.3925  ;
        POLYGON 0.0775 0.9775 0.8975 0.9775 0.8975 1.12 0.8325 1.12 0.8325 1.0425 0.1425 1.0425 0.1425 1.12 0.0775 1.12  ;
        POLYGON 0.0775 0.2775 0.1425 0.2775 0.1425 0.5225 0.8575 0.5225 0.8575 0.1925 1.2975 0.1925 1.2975 0.3625 1.2325 0.3625 1.2325 0.2575 0.9225 0.2575 0.9225 0.5875 0.0775 0.5875  ;
  END
END OAI222_X1

MACRO OAI222_X2
  CLASS core ;
  FOREIGN OAI222_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.52 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2625 1.315 0.2625 1.275 0.2625 1.045 0.3275 1.045 0.3275 1.275 0.3275 1.315 1.3625 1.315 1.3625 1.2475 1.3625 1.045 1.4275 1.045 1.4275 1.2475 1.4275 1.315 1.52 1.315 1.52 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.7025 0.6975 0.7025 0.7525 0.7025 0.7525 0.8375 0.6975 0.8375 0.6325 0.8375  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.8225 0.7025 0.8875 0.7025 1.0025 0.7025 1.0025 0.7625 1.0025 0.8375 0.9375 0.8375 0.8875 0.8375 0.8225 0.8375  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.2025 0.5625 1.2675 0.5625 1.2675 0.6975 1.2025 0.6975  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6125 1.045 0.6475 1.045 0.7125 1.045 0.7475 1.045 0.7475 1.185 0.9875 1.185 0.9875 0.9775 0.9875 0.9675 0.9875 0.9025 1.0725 0.9025 1.0725 0.51 1.0475 0.51 1.0475 0.3225 1.0725 0.3225 1.1125 0.3225 1.1125 0.4575 1.1375 0.4575 1.1375 0.8425 1.2675 0.8425 1.2675 0.9775 1.1375 0.9775 1.0725 0.9775 1.0525 0.9775 1.0525 1.25 0.7125 1.25 0.6475 1.25 0.6125 1.25 0.6125 1.11  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.7025 0.5075 0.7025 0.5625 0.7025 0.5625 0.8375 0.5075 0.8375 0.4425 0.8375  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4225 0.2625 0.4575 0.2625 0.4575 0.085 0 0.085 0 -0.085 1.52 -0.085 1.52 0.085 0.5225 0.085 0.5225 0.2625 0.5575 0.2625 0.5575 0.3275 0.5225 0.3275 0.4575 0.3275 0.4225 0.3275  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.7025 0.1275 0.7025 0.1275 0.8375 0.0625 0.8375  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.7025 0.3725 0.7025 0.3725 0.8375 0.2525 0.8375  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.2675 0.1825 0.3325 0.1825 0.3325 0.3925 0.6425 0.3925 0.6425 0.1825 0.7075 0.1825 0.7075 0.3925 0.7075 0.4275 0.7075 0.4575 0.2675 0.4575 0.2675 0.4275 0.2675 0.3925  ;
        POLYGON 0.0775 0.9025 0.8975 0.9025 0.8975 1.12 0.8325 1.12 0.8325 0.98 0.1425 0.98 0.1425 1.1775 0.0775 1.1775 0.0775 0.98 0.0775 0.965  ;
        POLYGON 0.0775 0.2025 0.1425 0.2025 0.1425 0.2375 0.1425 0.5225 0.8575 0.5225 0.8575 0.1925 1.2975 0.1925 1.2975 0.4775 1.2325 0.4775 1.2325 0.2575 0.9225 0.2575 0.9225 0.5875 0.0775 0.5875 0.0775 0.2375  ;
  END
END OAI222_X2

MACRO OAI222_X4
  CLASS core ;
  FOREIGN OAI222_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.66 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.0675 0.11 1.0675 0.11 1.315 0.765 1.315 0.765 1.2075 0.9 1.2075 0.9 1.315 1.56 1.315 1.56 1.0675 1.625 1.0675 1.625 1.315 2.08 1.315 2.08 1.1625 2.215 1.1625 2.215 1.315 2.66 1.315 2.66 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.0125 0.7975 1.2 0.7975 1.2 0.8425 1.2 0.8625 1.0775 0.8625 1.0775 0.9775 1.0125 0.9775 1.0125 0.8425  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.87 0.6225 2.51 0.6225 2.51 0.6875 2.4075 0.6875 2.4075 0.8375 2.3425 0.8375 2.3425 0.6875 1.87 0.6875  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.0825 0.7525 2.2525 0.7525 2.2525 0.8775 2.2525 0.9425 2.1175 0.9425 2.1175 0.8775 2.1175 0.8175 2.0825 0.8175  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.805 1.0325 2.46 1.0325 2.46 0.8775 2.595 0.8775 2.595 1.0975 1.705 1.0975 1.705 1.0025 1.485 1.0025 1.485 1.1425 0.39 1.1425 0.39 0.9275 0.525 0.9275 0.525 1.0775 1.42 1.0775 1.42 0.9375 1.74 0.9375 1.74 0.51 1.76 0.51 1.76 0.3775 1.725 0.3775 1.725 0.3125 1.86 0.3125 1.86 0.3775 1.825 0.3775 1.825 0.4925 2.1 0.4925 2.1 0.3125 2.235 0.3125 2.235 0.4925 2.515 0.4925 2.515 0.2775 2.58 0.2775 2.58 0.5575 1.805 0.5575  ;
    END
  END ZN
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.7975 0.415 0.7975 0.415 0.8625 0.1275 0.8625 0.1275 0.9775 0.0625 0.9775  ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.66 -0.085 2.66 0.085 0.675 0.085 0.675 0.425 0.61 0.425 0.61 0.085 0.295 0.085 0.295 0.425 0.23 0.425 0.23 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.875 0.6675 1.555 0.6675 1.555 0.7325 1.4575 0.7325 1.4575 0.8375 1.3925 0.8375 1.3925 0.7325 0.875 0.7325  ;
    END
  END B2
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.115 0.6675 0.795 0.6675 0.795 0.7325 0.6975 0.7325 0.6975 0.8375 0.6325 0.8375 0.6325 0.7325 0.115 0.7325  ;
    END
  END C2
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.2775 0.11 0.2775 0.11 0.49 0.42 0.49 0.42 0.2775 0.485 0.2775 0.485 0.49 0.8 0.49 0.8 0.2775 0.865 0.2775 0.865 0.49 1.145 0.49 1.145 0.3125 1.28 0.3125 1.28 0.49 1.525 0.49 1.525 0.3125 1.66 0.3125 1.66 0.5175 1.625 0.5175 1.625 0.555 0.09 0.555 0.09 0.5525 0.045 0.5525  ;
        POLYGON 0.995 0.15 2.39 0.15 2.39 0.425 2.325 0.425 2.325 0.215 2.01 0.215 2.01 0.425 1.945 0.425 1.945 0.215 1.435 0.215 1.435 0.425 1.37 0.425 1.37 0.215 1.06 0.215 1.06 0.425 0.995 0.425  ;
  END
END OAI222_X4

MACRO OAI22_X1
  CLASS core ;
  FOREIGN OAI22_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.14 0.11 1.14 0.11 1.315 0.8 1.315 0.8 1.14 0.865 1.14 0.865 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.5625 0.34 0.5625 0.34 0.6975 0.2525 0.6975  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.5625 0.53 0.5625 0.53 0.6975 0.4425 0.6975  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.295 0.085 0.295 0.3675 0.23 0.3675 0.23 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.8425 0.1275 0.8425 0.1275 0.9775 0.0625 0.9775  ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.5975 1.0175 0.695 1.0175 0.695 0.8925 0.8225 0.8925 0.8225 0.8425 0.8875 0.8425 0.8875 0.9575 0.76 0.9575 0.76 1.0825 0.5975 1.0825  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.425 0.7925 0.435 0.7925 0.435 0.7625 0.615 0.7625 0.615 0.2875 0.68 0.2875 0.68 0.5625 0.6975 0.5625 0.6975 0.6975 0.68 0.6975 0.68 0.8275 0.49 0.8275 0.49 1.1525 0.425 1.1525  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.2875 0.11 0.2875 0.11 0.4325 0.42 0.4325 0.42 0.1575 0.865 0.1575 0.865 0.3675 0.8 0.3675 0.8 0.2225 0.485 0.2225 0.485 0.4975 0.045 0.4975  ;
  END
END OAI22_X1

MACRO OAI22_X2
  CLASS core ;
  FOREIGN OAI22_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.0675 1.315 0.0675 1.0675 0.1325 1.0675 0.1325 1.315 0.8225 1.315 0.8225 1.0675 0.8875 1.0675 0.8875 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.5625 0.315 0.5625 0.3175 0.5625 0.4375 0.5625 0.4375 0.6375 0.3175 0.6375 0.3175 0.6975 0.2525 0.6975  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.7375 0.5025 0.7375 0.5025 0.6975 0.5675 0.6975 0.5675 0.7375 0.5675 0.8025 0.5675 0.8325 0.5025 0.8325 0.5025 0.8025 0.4075 0.8025  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.3175 0.085 0.3175 0.3625 0.2525 0.3625 0.2525 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1125 0.7975 0.2475 0.7975 0.2475 0.8775 0.3525 0.8775 0.3525 0.9425 0.1825 0.9425 0.1825 0.8625 0.1125 0.8625  ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.7625 0.7625 0.8225 0.7625 0.8225 0.7025 0.8875 0.7025 0.8875 0.8375 0.8275 0.8375 0.8275 0.8975 0.8225 0.8975 0.7625 0.8975  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 1.0175 0.4475 1.0175 0.4475 0.8975 0.6325 0.8975 0.6325 0.3725 0.5975 0.3725 0.5975 0.3075 0.7325 0.3075 0.7325 0.3725 0.6975 0.3725 0.6975 0.9625 0.5425 0.9625 0.5425 1.1375 0.4075 1.1375  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.0675 0.2725 0.1325 0.2725 0.1325 0.4275 0.4425 0.4275 0.4425 0.1775 0.8875 0.1775 0.8875 0.5025 0.8225 0.5025 0.8225 0.2425 0.5075 0.2425 0.5075 0.4925 0.0675 0.4925  ;
  END
END OAI22_X2

MACRO OAI22_X4
  CLASS core ;
  FOREIGN OAI22_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.9 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.1275 1.315 0.1275 1.0675 0.1925 1.0675 0.1925 1.315 0.8825 1.315 0.8825 1.0675 0.9475 1.0675 0.9475 1.315 1.6625 1.315 1.6625 1.0675 1.7275 1.0675 1.7275 1.315 1.9 1.315 1.9 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.8775 0.2875 0.8775 0.2875 0.7975 0.4575 0.7975 0.4575 0.8625 0.3525 0.8625 0.3525 0.9425 0.2175 0.9425  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.3325 0.7975 1.6475 0.7975 1.6475 0.9775 1.5825 0.9775 1.5825 0.8625 1.3325 0.8625  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.9 -0.085 1.9 0.085 0.7275 0.085 0.7275 0.4725 0.5925 0.4725 0.5925 0.085 0.3475 0.085 0.3475 0.4725 0.2125 0.4725 0.2125 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1725 0.6675 0.8025 0.6675 0.8025 0.8025 0.5975 0.8025 0.5975 0.7325 0.1725 0.7325  ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.0525 0.6675 1.6575 0.6675 1.6575 0.7325 1.2675 0.7325 1.2675 0.8375 1.2025 0.8375 1.2025 0.8025 1.0525 0.8025  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.5075 0.905 0.5975 0.905 0.5975 0.8775 0.9225 0.8775 0.9225 0.5375 1.035 0.5375 1.035 0.3125 1.17 0.3125 1.17 0.5375 1.435 0.5375 1.435 0.3125 1.57 0.3125 1.57 0.5625 1.495 0.5625 1.495 0.6025 0.9875 0.6025 0.9875 0.9275 1.3475 0.9275 1.3475 1.2025 1.2825 1.2025 1.2825 0.9925 0.5725 0.9925 0.5725 1.18 0.5075 1.18  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.0625 0.2775 0.1275 0.2775 0.1275 0.5375 0.4375 0.5375 0.4375 0.2775 0.5025 0.2775 0.5025 0.5375 0.7925 0.5375 0.7925 0.4175 0.8225 0.4175 0.8225 0.2675 0.8925 0.2675 0.8925 0.1825 1.72 0.1825 1.72 0.5075 1.655 0.5075 1.655 0.2475 1.37 0.2475 1.37 0.4725 1.235 0.4725 1.235 0.2475 0.9575 0.2475 0.9575 0.4725 0.8575 0.4725 0.8575 0.5975 0.8175 0.5975 0.8175 0.6025 0.0625 0.6025  ;
  END
END OAI22_X4

MACRO OAI33_X1
  CLASS core ;
  FOREIGN OAI33_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.085 1.315 0.085 0.995 0.15 0.995 0.15 1.315 1.22 1.315 1.22 0.995 1.285 0.995 1.285 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.5975 0.595 0.5975 0.595 0.7325 0.53 0.7325 0.53 0.6625 0.4075 0.6625  ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.785 0.825 0.85 0.825 0.85 1.1575 0.9225 1.1575 0.9225 1.2225 0.785 1.2225  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.95 0.5975 1.1125 0.5975 1.1125 0.6625 1.015 0.6625 1.015 0.7325 0.95 0.7325  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.655 0.775 0.66 0.775 0.66 0.61 0.675 0.61 0.675 0.5875 0.82 0.5875 0.82 0.475 0.84 0.475 0.84 0.3125 0.905 0.3125 0.905 0.4575 1.22 0.4575 1.22 0.3125 1.285 0.3125 1.285 0.5225 0.885 0.5225 0.885 0.6525 0.725 0.6525 0.725 0.8 0.72 0.8 0.72 1.225 0.655 1.225  ;
    END
  END ZN
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.9775 0.8775 1.115 0.8775 1.115 0.8075 1.18 0.8075 1.18 0.9425 0.9775 0.9425  ;
    END
  END A3
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.5975 0.1625 0.5975 0.1625 0.6625 0.1275 0.6625 0.1275 0.8375 0.0625 0.8375  ;
    END
  END B3
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 0.525 0.085 0.525 0.3925 0.46 0.3925 0.46 0.085 0.15 0.085 0.15 0.3925 0.085 0.3925 0.085 0.085 0 0.085  ;
    END
  END VSS
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.355 0.825 0.5075 0.825 0.5075 0.9775 0.355 0.9775  ;
    END
  END B2
  OBS
      LAYER metal1 ;
        POLYGON 0.275 0.3125 0.34 0.3125 0.34 0.4575 0.65 0.4575 0.65 0.1825 1.095 0.1825 1.095 0.3925 1.03 0.3925 1.03 0.2475 0.715 0.2475 0.715 0.5225 0.275 0.5225  ;
  END
END OAI33_X1

MACRO OR2_X1
  CLASS core ;
  FOREIGN OR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.46 1.315 0.46 1.115 0.525 1.115 0.525 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.215 0.7375 0.3525 0.7375 0.3525 0.8025 0.28 0.8025 0.28 0.8725 0.215 0.8725  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.525 0.085 0.525 0.3325 0.46 0.3325 0.46 0.085 0.15 0.085 0.15 0.3325 0.085 0.3325 0.085 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.355 0.8675 0.5425 0.8675 0.5425 0.9425 0.42 0.9425 0.42 1.0025 0.355 1.0025  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.5975 0.65 0.5975 0.65 0.2125 0.715 0.2125 0.715 1.19 0.65 1.19 0.65 0.6625 0.4075 0.6625  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.085 0.42 0.1 0.42 0.1 0.3975 0.27 0.3975 0.27 0.2125 0.335 0.2125 0.335 0.3975 0.585 0.3975 0.585 0.5325 0.52 0.5325 0.52 0.4625 0.15 0.4625 0.15 1.1275 0.085 1.1275  ;
  END
END OR2_X1

MACRO OR2_X2
  CLASS core ;
  FOREIGN OR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.4475 1.315 0.4475 0.99 0.5125 0.99 0.5125 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1825 0.5275 0.2475 0.5275 0.2475 0.5975 0.5425 0.5975 0.5425 0.6625 0.1825 0.6625  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.5075 0.085 0.5075 0.3325 0.4425 0.3325 0.4425 0.085 0.1325 0.085 0.1325 0.3325 0.0675 0.3325 0.0675 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.8775 0.3375 0.8775 0.3375 0.8075 0.4025 0.8075 0.4025 0.9425 0.2175 0.9425  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.2725 0.6975 0.2725 0.6975 1.21 0.6325 1.21  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.0525 0.3975 0.2525 0.3975 0.2525 0.2125 0.3175 0.2125 0.3175 0.3975 0.5675 0.3975 0.5675 0.5325 0.5025 0.5325 0.5025 0.4625 0.1175 0.4625 0.1175 1.1425 0.0525 1.1425  ;
  END
END OR2_X2

MACRO OR2_X4
  CLASS core ;
  FOREIGN OR2_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.4475 1.315 0.4475 1.0075 0.5125 1.0075 0.5125 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1825 0.9 0.2475 0.9 0.2475 1.1575 0.3525 1.1575 0.3525 1.2225 0.1825 1.2225  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.5125 0.085 0.5125 0.4075 0.4475 0.4075 0.4475 0.085 0.1175 0.085 0.1175 0.5375 0.0525 0.5375 0.0525 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3225 0.7875 0.3875 0.7875 0.3875 0.8775 0.5425 0.8775 0.5425 0.9425 0.3225 0.9425  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.2775 0.6975 0.2775 0.6975 0.9575 0.6325 0.9575  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.0525 0.635 0.0675 0.635 0.0675 0.6125 0.2375 0.6125 0.2375 0.4175 0.3025 0.4175 0.3025 0.6125 0.5025 0.6125 0.5025 0.5425 0.5675 0.5425 0.5675 0.6775 0.1175 0.6775 0.1175 1.16 0.0525 1.16  ;
  END
END OR2_X4

MACRO OR3_X1
  CLASS core ;
  FOREIGN OR3_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.6175 1.315 0.6175 1.0025 0.6825 1.0025 0.6825 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.8775 0.5275 0.8775 0.5275 0.8075 0.5925 0.8075 0.5925 0.9425 0.4075 0.9425  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1825 0.6675 0.2475 0.6675 0.2475 0.7375 0.3525 0.7375 0.3525 0.8025 0.1825 0.8025  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.6975 0.085 0.6975 0.3425 0.6325 0.3425 0.6325 0.085 0.3175 0.085 0.3175 0.3425 0.2525 0.3425 0.2525 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3375 0.5375 0.4025 0.5375 0.4025 0.5975 0.5425 0.5975 0.5425 0.6725 0.3375 0.6725  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.8225 0.2225 0.8875 0.2225 0.8875 1.2175 0.8225 1.2175  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.0525 0.43 0.0675 0.43 0.0675 0.2225 0.1325 0.2225 0.1325 0.4075 0.4425 0.4075 0.4425 0.2225 0.5075 0.2225 0.5075 0.4075 0.7575 0.4075 0.7575 0.5425 0.6925 0.5425 0.6925 0.4725 0.1175 0.4725 0.1175 1.2325 0.0525 1.2325  ;
  END
END OR3_X1

MACRO OR3_X2
  CLASS core ;
  FOREIGN OR3_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.61 1.315 0.61 0.995 0.675 0.995 0.675 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.8775 0.505 0.8775 0.505 0.8075 0.57 0.8075 0.57 0.9425 0.4075 0.9425  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.6675 0.24 0.6675 0.24 0.7375 0.3525 0.7375 0.3525 0.8025 0.175 0.8025  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.675 0.085 0.675 0.2975 0.61 0.2975 0.61 0.085 0.295 0.085 0.295 0.2975 0.23 0.2975 0.23 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.34 0.5275 0.405 0.5275 0.405 0.5975 0.5425 0.5975 0.5425 0.6625 0.34 0.6625  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.5625 0.8 0.5625 0.8 0.2375 0.865 0.2375 0.865 1.215 0.8 1.215 0.8 0.6975 0.6325 0.6975  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.1775 0.11 0.1775 0.11 0.3625 0.42 0.3625 0.42 0.1775 0.485 0.1775 0.485 0.3625 0.735 0.3625 0.735 0.4975 0.67 0.4975 0.67 0.4275 0.11 0.4275 0.11 1.225 0.045 1.225  ;
  END
END OR3_X2

MACRO OR3_X4
  CLASS core ;
  FOREIGN OR3_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.95 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.625 1.315 0.625 0.9375 0.69 0.9375 0.69 1.315 0.95 1.315 0.95 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4425 0.5625 0.53 0.5625 0.53 0.6975 0.4425 0.6975  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.19 0.5625 0.3175 0.5625 0.3175 0.6975 0.19 0.6975  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.95 -0.085 0.95 0.085 0.695 0.085 0.695 0.3525 0.63 0.3525 0.63 0.085 0.295 0.085 0.295 0.3675 0.23 0.3675 0.23 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.7675 0.355 0.7675 0.355 0.9775 0.2525 0.9775  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.815 0.2225 0.88 0.2225 0.88 0.5625 0.8875 0.5625 0.8875 0.6975 0.88 0.6975 0.88 0.8875 0.815 0.8875  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.2475 0.11 0.2475 0.11 0.4325 0.42 0.4325 0.42 0.2475 0.485 0.2475 0.485 0.4325 0.75 0.4325 0.75 0.6225 0.685 0.6225 0.685 0.4975 0.125 0.4975 0.125 1.1675 0.06 1.1675 0.06 0.475 0.045 0.475  ;
  END
END OR3_X4

MACRO OR4_X1
  CLASS core ;
  FOREIGN OR4_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.8075 1.315 0.8075 0.9375 0.8725 0.9375 0.8725 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4975 0.5975 0.7325 0.5975 0.7325 0.6625 0.4975 0.6625  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1825 0.5625 0.2475 0.5625 0.2475 0.5975 0.3525 0.5975 0.3525 0.6625 0.2475 0.6625 0.2475 0.6975 0.1825 0.6975  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.8875 0.085 0.8875 0.3525 0.8225 0.3525 0.8225 0.085 0.5075 0.085 0.5075 0.3525 0.4425 0.3525 0.4425 0.085 0.1325 0.085 0.1325 0.3525 0.0675 0.3525 0.0675 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3025 0.7375 0.5425 0.7375 0.5425 0.8025 0.3025 0.8025  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6825 0.7375 0.9225 0.7375 0.9225 0.8025 0.6825 0.8025  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.0125 0.2325 1.0775 0.2325 1.0775 1.1525 1.0125 1.1525  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.0525 0.4175 0.2525 0.4175 0.2525 0.2325 0.3175 0.2325 0.3175 0.4175 0.6325 0.4175 0.6325 0.2325 0.6975 0.2325 0.6975 0.4175 0.9475 0.4175 0.9475 0.5525 0.8825 0.5525 0.8825 0.4825 0.1175 0.4825 0.1175 1.1025 0.0525 1.1025  ;
  END
END OR4_X1

MACRO OR4_X2
  CLASS core ;
  FOREIGN OR4_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.8075 1.315 0.8075 0.9375 0.8725 0.9375 0.8725 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4975 0.5975 0.7325 0.5975 0.7325 0.6625 0.4975 0.6625  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1825 0.5625 0.2475 0.5625 0.2475 0.5975 0.3525 0.5975 0.3525 0.6625 0.2475 0.6625 0.2475 0.6975 0.1825 0.6975  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.8875 0.085 0.8875 0.3525 0.8225 0.3525 0.8225 0.085 0.5075 0.085 0.5075 0.3525 0.4425 0.3525 0.4425 0.085 0.1325 0.085 0.1325 0.3525 0.0675 0.3525 0.0675 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3025 0.7375 0.5425 0.7375 0.5425 0.8025 0.3025 0.8025  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6825 0.7375 0.9225 0.7375 0.9225 0.8025 0.6825 0.8025  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.0125 0.2325 1.0775 0.2325 1.0775 1.0175 1.0125 1.0175  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.0525 0.4175 0.2525 0.4175 0.2525 0.2325 0.3175 0.2325 0.3175 0.4175 0.6325 0.4175 0.6325 0.2325 0.6975 0.2325 0.6975 0.4175 0.9475 0.4175 0.9475 0.5525 0.8825 0.5525 0.8825 0.4825 0.1175 0.4825 0.1175 1.1025 0.0525 1.1025  ;
  END
END OR4_X2

MACRO OR4_X4
  CLASS core ;
  FOREIGN OR4_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.8075 1.315 0.8075 0.9375 0.8725 0.9375 0.8725 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4975 0.5975 0.7325 0.5975 0.7325 0.6625 0.4975 0.6625  ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1825 0.5625 0.2475 0.5625 0.2475 0.5975 0.3525 0.5975 0.3525 0.6625 0.2475 0.6625 0.2475 0.6975 0.1825 0.6975  ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.8875 0.085 0.8875 0.3525 0.8225 0.3525 0.8225 0.085 0.5075 0.085 0.5075 0.3525 0.4425 0.3525 0.4425 0.085 0.1325 0.085 0.1325 0.3525 0.0675 0.3525 0.0675 0.085 0 0.085  ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3025 0.7375 0.5425 0.7375 0.5425 0.8025 0.3025 0.8025  ;
    END
  END A2
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6825 0.7375 0.9225 0.7375 0.9225 0.8025 0.6825 0.8025  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.0125 0.165 1.0775 0.165 1.0775 1.1675 1.0125 1.1675  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.0525 0.4175 0.2525 0.4175 0.2525 0.2325 0.3175 0.2325 0.3175 0.4175 0.6325 0.4175 0.6325 0.2325 0.6975 0.2325 0.6975 0.4175 0.9475 0.4175 0.9475 0.565 0.8825 0.565 0.8825 0.4825 0.1175 0.4825 0.1175 1.1025 0.0525 1.1025  ;
  END
END OR4_X4

MACRO SDFFRS_X1
  CLASS core ;
  FOREIGN SDFFRS_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 6.65 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 5.9175 0.37 6.0525 0.37 6.0525 0.7125 5.9175 0.7125  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.1025 0.5675 3.2575 0.5675 3.2575 0.4575 3.3925 0.4575 3.3925 0.57 5.0225 0.57 5.0225 0.635 3.3725 0.635 3.3725 0.6325 3.1025 0.6325  ;
    END
  END SN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1775 1.0175 0.3525 1.0175 0.3525 1.0825 0.1775 1.0825  ;
    END
  END SE
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.6975 0.71 4.895 0.71 4.895 0.775 3.6975 0.775  ;
        POLYGON 5.4825 0.9025 5.8725 0.9025 5.8725 0.9675 5.43 0.9675 5.43 0.9425 5.3475 0.9425 5.3475 0.7375 5.4175 0.7375 5.4175 0.4625 5.5525 0.4625 5.5525 0.5275 5.4825 0.5275  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 6.3125 1.315 6.65 1.315 6.65 1.485 0 1.485 0 1.315 0.3025 1.315 0.3025 1.1475 0.4375 1.1475 0.4375 1.315 1.0575 1.315 1.0575 1.1475 1.1925 1.1475 1.1925 1.315 1.62 1.315 1.62 1.1075 1.755 1.1075 1.755 1.315 2.4325 1.315 2.4325 1.175 2.3625 1.175 2.3625 1.11 2.4975 1.11 2.4975 1.315 3.3975 1.315 3.3975 1.175 3.3275 1.175 3.3275 1.11 3.4625 1.11 3.4625 1.315 3.8475 1.315 3.8475 1.175 3.7775 1.175 3.7775 1.11 3.9125 1.11 3.9125 1.315 4.53 1.315 4.53 1.1925 4.665 1.1925 4.665 1.315 5.3875 1.315 5.3875 1.1925 5.5225 1.1925 5.5225 1.315 5.8175 1.315 5.8175 1.1925 5.9525 1.1925 5.9525 1.315 6.2475 1.315 6.2475 0.7075 6.3825 0.7075 6.3825 0.7725 6.3125 0.7725  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 6.4475 0.6475 6.5225 0.6475 6.5225 0.435 6.4475 0.435 6.4475 0.37 6.5875 0.37 6.5875 0.7125 6.4475 0.7125  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.3175 0.5425 0.3175 0.5425 0.385 0.9875 0.385 0.9875 0.645 0.9225 0.645 0.9225 0.45 0.4075 0.45  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 6.65 -0.085 6.65 0.085 6.3825 0.085 6.3825 0.42 6.2475 0.42 6.2475 0.085 5.3775 0.085 5.3775 0.1775 5.2425 0.1775 5.2425 0.085 4.9775 0.085 4.9775 0.235 4.8425 0.235 4.8425 0.085 3.9125 0.085 3.9125 0.235 3.7775 0.235 3.7775 0.085 3.1425 0.085 3.1425 0.2225 3.0075 0.2225 3.0075 0.085 2.1475 0.085 2.1475 0.2225 2.0125 0.2225 2.0125 0.085 1.765 0.085 1.765 0.2575 1.63 0.2575 1.63 0.085 1.235 0.085 1.235 0.19 1.1 0.19 1.1 0.085 0.4375 0.085 0.4375 0.19 0.3025 0.19 0.3025 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.71 1.055 0.71 1.055 0.385 1.12 0.385 1.12 0.775 0.5425 0.775 0.5425 0.8025 0.4075 0.8025  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.5475 0.4575 1.6825 0.4575 1.6825 0.5225 1.5475 0.5225  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.0975 0.8625 0.1675 0.8625 0.1675 0.215 0.0975 0.215 0.0975 0.15 0.2325 0.15 0.2325 0.515 0.8575 0.515 0.8575 0.58 0.2325 0.58 0.2325 0.9275 0.0975 0.9275  ;
        POLYGON 1.295 0.97 1.57 0.97 1.57 1.035 1.295 1.035  ;
        POLYGON 1.825 0.97 2.1 0.97 2.1 1.035 1.825 1.035  ;
        POLYGON 0.6825 0.8625 0.7925 0.8625 0.7925 0.84 1.185 0.84 1.185 0.32 0.8075 0.32 0.8075 0.295 0.725 0.295 0.725 0.23 0.86 0.23 0.86 0.255 1.25 0.255 1.25 0.84 2.2275 0.84 2.2275 0.905 0.8425 0.905 0.8425 0.9225 0.8175 0.9225 0.8175 0.9275 0.6825 0.9275  ;
        POLYGON 2.4325 0.5675 2.4925 0.5675 2.4925 0.4925 2.4225 0.4925 2.4225 0.4275 2.5575 0.4275 2.5575 0.5675 2.5675 0.5675 2.5675 0.6325 2.4325 0.6325  ;
        POLYGON 1.4825 0.6975 2.4175 0.6975 2.4175 0.825 2.8575 0.825 2.8575 0.89 2.3525 0.89 2.3525 0.7625 1.39 0.7625 1.39 0.6975 1.4175 0.6975 1.4175 0.2975 1.5775 0.2975 1.5775 0.3625 1.4825 0.3625  ;
        POLYGON 3.2125 0.1825 3.4875 0.1825 3.4875 0.2475 3.2125 0.2475  ;
        POLYGON 2.9775 0.7 3.3875 0.7 3.3875 0.7025 3.4325 0.7025 3.4325 0.84 3.6925 0.84 3.6925 0.905 3.3675 0.905 3.3675 0.765 2.9775 0.765  ;
        POLYGON 1.9875 1.11 2.2325 1.11 2.2325 0.98 2.4075 0.98 2.4075 0.97 2.5425 0.97 2.5425 0.98 2.9275 0.98 2.9275 0.97 4.3425 0.97 4.3425 1.035 2.9625 1.035 2.9625 1.16 2.8275 1.16 2.8275 1.045 2.2975 1.045 2.2975 1.175 1.9875 1.175  ;
        POLYGON 4.1825 0.185 4.3375 0.185 4.3375 0.31 4.5475 0.31 4.5475 0.375 4.2725 0.375 4.2725 0.25 4.1825 0.25  ;
        POLYGON 5.0175 0.8625 5.0875 0.8625 5.0875 0.505 4.1425 0.505 4.1425 0.38 2.6375 0.38 2.6375 0.3625 2.075 0.3625 2.075 0.4775 1.94 0.4775 1.94 0.3625 1.8175 0.3625 1.8175 0.2975 2.6825 0.2975 2.6825 0.315 4.2075 0.315 4.2075 0.44 5.1525 0.44 5.1525 0.9275 5.0175 0.9275  ;
        POLYGON 5.6825 0.7725 5.7475 0.7725 5.7475 0.8375 5.6125 0.8375 5.6125 0.7725 5.6175 0.7725 5.6175 0.3875 5.1925 0.3875 5.1925 0.375 4.6125 0.375 4.6125 0.31 5.2325 0.31 5.2325 0.3225 5.6925 0.3225 5.6925 0.3875 5.6825 0.3875  ;
        POLYGON 5.2825 1.0525 5.8725 1.0525 5.8725 1.1175 5.0875 1.1175 5.0875 1.2425 4.9525 1.2425 4.9525 1.1275 4.465 1.1275 4.465 1.1975 3.9775 1.1975 3.9775 1.1325 4.4 1.1325 4.4 1.0675 4.44 1.0675 4.44 1.0525 4.5775 1.0525 4.5775 1.0625 5.0525 1.0625 5.0525 1.0525 5.2175 1.0525 5.2175 0.4625 5.3525 0.4625 5.3525 0.5275 5.2825 0.5275  ;
        POLYGON 6.0275 1.1325 6.1175 1.1325 6.1175 0.2325 5.6375 0.2325 5.6375 0.1675 6.1825 0.1675 6.1825 0.5225 6.4225 0.5225 6.4225 0.5875 6.1825 0.5875 6.1825 1.1975 6.0275 1.1975  ;
  END
END SDFFRS_X1

MACRO SDFFRS_X2
  CLASS core ;
  FOREIGN SDFFRS_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 6.65 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 5.8675 0.6475 5.9375 0.6475 5.9375 0.3825 5.7275 0.3825 5.7275 0.3175 6.0025 0.3175 6.0025 0.7125 5.8675 0.7125  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.0325 0.55 3.2575 0.55 3.2575 0.4575 3.3925 0.4575 3.3925 0.555 4.9525 0.555 4.9525 0.62 3.3725 0.62 3.3725 0.6175 3.0325 0.6175  ;
    END
  END SN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1775 1.0175 0.3525 1.0175 0.3525 1.0825 0.1775 1.0825  ;
    END
  END SE
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.6275 0.6925 4.825 0.6925 4.825 0.7575 3.6275 0.7575  ;
        POLYGON 5.4125 0.8775 5.9325 0.8775 5.9325 0.9675 6.0025 0.9675 6.0025 1.0325 5.8675 1.0325 5.8675 0.9425 5.3475 0.9425 5.3475 0.785 5.2775 0.785 5.2775 0.72 5.3475 0.72 5.3475 0.445 5.4825 0.445 5.4825 0.51 5.4125 0.51  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 6.2625 1.315 6.65 1.315 6.65 1.485 0 1.485 0 1.315 0.3025 1.315 0.3025 1.1475 0.4375 1.1475 0.4375 1.315 1.0575 1.315 1.0575 1.1475 1.1925 1.1475 1.1925 1.315 1.55 1.315 1.55 1.09 1.685 1.09 1.685 1.315 2.3625 1.315 2.3625 1.1575 2.2925 1.1575 2.2925 1.0925 2.4275 1.0925 2.4275 1.315 3.3275 1.315 3.3275 1.1575 3.2575 1.1575 3.2575 1.0925 3.3925 1.0925 3.3925 1.315 3.7775 1.315 3.7775 1.1575 3.7075 1.1575 3.7075 1.0925 3.8425 1.0925 3.8425 1.315 4.46 1.315 4.46 1.175 4.595 1.175 4.595 1.315 5.3175 1.315 5.3175 1.175 5.4525 1.175 5.4525 1.315 5.7475 1.315 5.7475 1.175 5.8825 1.175 5.8825 1.315 6.1975 1.315 6.1975 0.8425 6.3325 0.8425 6.3325 0.9075 6.2625 0.9075  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 6.3825 0.6475 6.455 0.6475 6.455 0.4175 6.385 0.4175 6.385 0.3525 6.52 0.3525 6.52 0.4225 6.5875 0.4225 6.5875 0.5575 6.52 0.5575 6.52 0.7125 6.3825 0.7125  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.3175 0.5425 0.3175 0.5425 0.3675 0.9875 0.3675 0.9875 0.6275 0.9225 0.6275 0.9225 0.4325 0.4075 0.4325  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 6.1975 0.2475 6.2675 0.2475 6.2675 0.085 5.3075 0.085 5.3075 0.16 5.1725 0.16 5.1725 0.085 4.9075 0.085 4.9075 0.22 4.7725 0.22 4.7725 0.085 3.8425 0.085 3.8425 0.22 3.7075 0.22 3.7075 0.085 3.0725 0.085 3.0725 0.205 2.9375 0.205 2.9375 0.085 2.0775 0.085 2.0775 0.205 1.9425 0.205 1.9425 0.085 1.6975 0.085 1.6975 0.24 1.5625 0.24 1.5625 0.085 1.235 0.085 1.235 0.1725 1.1 0.1725 1.1 0.085 0.4375 0.085 0.4375 0.1725 0.3025 0.1725 0.3025 0.085 0 0.085 0 -0.085 6.65 -0.085 6.65 0.085 6.3325 0.085 6.3325 0.3125 6.1975 0.3125  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.6925 1.055 0.6925 1.055 0.3675 1.12 0.3675 1.12 0.7575 0.5425 0.7575 0.5425 0.8025 0.4075 0.8025  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.505 0.4575 1.6825 0.4575 1.6825 0.5225 1.505 0.5225  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.0975 0.8625 0.1675 0.8625 0.1675 0.215 0.0975 0.215 0.0975 0.15 0.2325 0.15 0.2325 0.4975 0.8575 0.4975 0.8575 0.5625 0.2325 0.5625 0.2325 0.9275 0.0975 0.9275  ;
        POLYGON 1.225 0.9525 1.5 0.9525 1.5 1.0175 1.225 1.0175  ;
        POLYGON 1.755 0.9525 2.03 0.9525 2.03 1.0175 1.755 1.0175  ;
        POLYGON 0.6825 0.8525 0.7925 0.8525 0.7925 0.8225 1.185 0.8225 1.185 0.3025 0.8075 0.3025 0.8075 0.2775 0.725 0.2775 0.725 0.2125 0.86 0.2125 0.86 0.2375 1.25 0.2375 1.25 0.8225 2.1575 0.8225 2.1575 0.8875 0.8475 0.8875 0.8475 0.9125 0.8175 0.9125 0.8175 0.9275 0.6825 0.9275  ;
        POLYGON 2.3625 0.55 2.4075 0.55 2.4075 0.475 2.3375 0.475 2.3375 0.41 2.4725 0.41 2.4725 0.55 2.4975 0.55 2.4975 0.615 2.3625 0.615  ;
        POLYGON 1.44 0.68 2.3475 0.68 2.3475 0.8075 2.7875 0.8075 2.7875 0.8725 2.2825 0.8725 2.2825 0.745 1.32 0.745 1.32 0.68 1.375 0.68 1.375 0.28 1.51 0.28 1.51 0.345 1.44 0.345  ;
        POLYGON 3.1425 0.165 3.4175 0.165 3.4175 0.23 3.1425 0.23  ;
        POLYGON 2.9075 0.6825 3.3175 0.6825 3.3175 0.685 3.3625 0.685 3.3625 0.8225 3.6225 0.8225 3.6225 0.8875 3.2975 0.8875 3.2975 0.7475 2.9075 0.7475  ;
        POLYGON 1.9175 1.0925 2.1625 1.0925 2.1625 0.9625 2.3375 0.9625 2.3375 0.9525 2.4725 0.9525 2.4725 0.9625 2.8575 0.9625 2.8575 0.9525 4.2725 0.9525 4.2725 1.0175 2.8925 1.0175 2.8925 1.1425 2.7575 1.1425 2.7575 1.0275 2.2275 1.0275 2.2275 1.1575 1.9175 1.1575  ;
        POLYGON 4.1125 0.1675 4.2675 0.1675 4.2675 0.295 4.4775 0.295 4.4775 0.36 4.2025 0.36 4.2025 0.2325 4.1125 0.2325  ;
        POLYGON 4.9475 0.845 5.0175 0.845 5.0175 0.49 4.0725 0.49 4.0725 0.3625 2.5675 0.3625 2.5675 0.345 2.005 0.345 2.005 0.4625 1.87 0.4625 1.87 0.345 1.75 0.345 1.75 0.28 2.6125 0.28 2.6125 0.2975 4.1375 0.2975 4.1375 0.425 5.0825 0.425 5.0825 0.91 4.9475 0.91  ;
        POLYGON 5.6125 0.7475 5.6625 0.7475 5.6625 0.8125 5.5275 0.8125 5.5275 0.7475 5.5475 0.7475 5.5475 0.37 5.1175 0.37 5.1175 0.36 4.5425 0.36 4.5425 0.295 5.1525 0.295 5.1525 0.305 5.6225 0.305 5.6225 0.37 5.6125 0.37  ;
        POLYGON 5.2125 1.035 5.8025 1.035 5.8025 1.1 4.9975 1.1 4.9975 1.225 4.8625 1.225 4.8625 1.11 4.395 1.11 4.395 1.18 3.9075 1.18 3.9075 1.115 4.33 1.115 4.33 1.05 4.37 1.05 4.37 1.035 4.5075 1.035 4.5075 1.045 4.9625 1.045 4.9625 1.035 5.1475 1.035 5.1475 0.445 5.2825 0.445 5.2825 0.51 5.2125 0.51  ;
        POLYGON 5.9775 1.115 6.0675 1.115 6.0675 0.215 5.5675 0.215 5.5675 0.15 6.1325 0.15 6.1325 0.48 6.365 0.48 6.365 0.545 6.1325 0.545 6.1325 1.18 5.9775 1.18  ;
  END
END SDFFRS_X2

MACRO SDFFR_X1
  CLASS core ;
  FOREIGN SDFFR_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 4.94 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.15 0.1275 0.15 0.1275 1.2375 0.0625 1.2375  ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 4.6225 0.6575 4.6875 0.6575 4.6875 0.8375 4.6225 0.8375  ;
    END
  END SE
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.3925 0.7025 1.4575 0.7025 1.4575 0.85 2.6325 0.85 2.6325 0.915 1.3925 0.915  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2475 1.315 0.2475 1.0175 0.3125 1.0175 0.3125 1.315 0.7775 1.315 0.7775 1.13 0.8425 1.13 0.8425 1.315 1.5025 1.315 1.5025 1.2425 1.6375 1.2425 1.6375 1.315 2.2575 1.315 2.2575 1.13 2.3225 1.13 2.3225 1.315 2.6725 1.315 2.6725 1.19 2.6025 1.19 2.6025 1.125 2.7375 1.125 2.7375 1.315 3.4175 1.315 3.4175 1.09 3.4825 1.09 3.4825 1.185 3.8075 1.185 3.8075 1.1025 3.9425 1.1025 3.9425 1.315 4.5975 1.315 4.5975 1.0675 4.6625 1.0675 4.6625 1.315 4.94 1.315 4.94 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.7025 0.4375 0.7025 0.4375 0.15 0.5025 0.15 0.5025 1.2375 0.4375 1.2375 0.4375 0.8375 0.2525 0.8375  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.9525 0.5425 4.57 0.5425 4.57 0.6075 4.1175 0.6075 4.1175 0.6975 4.0525 0.6975 4.0525 0.6425 3.9525 0.6425  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 4.94 -0.085 4.94 0.085 4.64 0.085 4.64 0.1925 4.575 0.1925 4.575 0.085 3.8225 0.085 3.8225 0.1925 3.7575 0.1925 3.7575 0.085 3.4775 0.085 3.4775 0.1925 3.4125 0.1925 3.4125 0.085 2.7525 0.085 2.7525 0.235 2.6175 0.235 2.6175 0.085 1.8825 0.085 1.8825 0.1925 1.8175 0.1925 1.8175 0.085 0.9175 0.085 0.9175 0.27 0.8525 0.27 0.8525 0.085 0.3125 0.085 0.3125 0.27 0.2475 0.27 0.2475 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.8625 0.7025 3.9275 0.7025 3.9275 0.8425 4.4125 0.8425 4.4125 0.9225 4.5925 0.9225 4.5925 0.9875 4.3475 0.9875 4.3475 0.9075 3.8625 0.9075  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.4825 0.7025 3.5475 0.7025 3.5475 0.8375 3.4825 0.8375  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.5725 0.3725 0.6475 0.3725 0.6475 0.1625 0.7125 0.1625 0.7125 0.4375 0.6375 0.4375 0.6375 1.115 0.6575 1.115 0.6575 1.25 0.5725 1.25  ;
        POLYGON 1.17 1.1125 1.9825 1.1125 1.9825 1.2475 1.9175 1.2475 1.9175 1.1775 1.2225 1.1775 1.2225 1.25 1.1575 1.25 1.1575 1.1775 1.105 1.1775 1.105 0.5275 0.8375 0.5275 0.8375 0.8025 0.7025 0.8025 0.7025 0.7375 0.7725 0.7375 0.7725 0.4625 1.105 0.4625 1.105 0.22 1.4175 0.22 1.4175 0.15 1.4825 0.15 1.4825 0.285 1.17 0.285  ;
        POLYGON 2.2775 0.15 2.3425 0.15 2.3425 0.31 2.8125 0.31 2.8125 0.375 2.2775 0.375  ;
        POLYGON 2.4525 0.9925 2.4775 0.9925 2.4775 0.98 2.8125 0.98 2.8125 1.045 2.5175 1.045 2.5175 1.25 2.4525 1.25  ;
        POLYGON 1.235 0.35 2.0025 0.35 2.0025 0.1625 2.0675 0.1625 2.0675 0.44 2.9675 0.44 2.9675 0.505 2.0025 0.505 2.0025 0.415 1.3 0.415 1.3 0.9825 2.1375 0.9825 2.1375 1.2375 2.0725 1.2375 2.0725 1.0475 1.235 1.0475  ;
        POLYGON 1.7125 0.5725 3.0325 0.5725 3.0325 0.15 3.0975 0.15 3.0975 0.6125 3.1025 0.6125 3.1025 1.12 3.0375 1.12 3.0375 0.6375 1.7125 0.6375  ;
        POLYGON 3.2325 0.96 3.6675 0.96 3.6675 1.12 3.6025 1.12 3.6025 1.025 3.2325 1.025 3.2325 1.25 2.9075 1.25 2.9075 0.92 2.8375 0.92 2.8375 0.785 1.5825 0.785 1.5825 0.545 1.365 0.545 1.365 0.48 1.6475 0.48 1.6475 0.72 2.9025 0.72 2.9025 0.855 2.9725 0.855 2.9725 1.185 3.1675 1.185 3.1675 0.2575 3.6025 0.2575 3.6025 0.1625 3.6675 0.1625 3.6675 0.3225 3.2325 0.3225  ;
        POLYGON 3.7975 0.9725 4.2825 0.9725 4.2825 1.1475 4.2175 1.1475 4.2175 1.0375 3.7325 1.0375 3.7325 0.6375 3.2975 0.6375 3.2975 0.5725 3.7325 0.5725 3.7325 0.3225 3.7375 0.3225 3.7375 0.2825 4.1925 0.2825 4.1925 0.1625 4.2575 0.1625 4.2575 0.3475 3.7975 0.3475  ;
        POLYGON 4.0775 0.4125 4.765 0.4125 4.765 0.1625 4.83 0.1625 4.83 0.4275 4.8525 0.4275 4.8525 1.1475 4.7875 1.1475 4.7875 0.4775 4.0775 0.4775  ;
  END
END SDFFR_X1

MACRO SDFFR_X2
  CLASS core ;
  FOREIGN SDFFR_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 4.94 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.2125 0.1275 0.2125 0.1275 1.2375 0.0625 1.2375  ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 4.6225 0.6575 4.6875 0.6575 4.6875 0.8375 4.6225 0.8375  ;
    END
  END SE
  PIN RN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.3925 0.7025 1.4575 0.7025 1.4575 0.85 2.6325 0.85 2.6325 0.915 1.3925 0.915  ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2475 1.315 0.2475 1.0175 0.3125 1.0175 0.3125 1.315 0.7775 1.315 0.7775 1.13 0.8425 1.13 0.8425 1.315 1.5025 1.315 1.5025 1.2425 1.6375 1.2425 1.6375 1.315 2.2575 1.315 2.2575 1.13 2.3225 1.13 2.3225 1.315 2.6725 1.315 2.6725 1.19 2.6025 1.19 2.6025 1.125 2.7375 1.125 2.7375 1.315 3.4175 1.315 3.4175 1.09 3.4825 1.09 3.4825 1.185 3.8075 1.185 3.8075 1.1025 3.9425 1.1025 3.9425 1.315 4.5975 1.315 4.5975 1.0675 4.6625 1.0675 4.6625 1.315 4.94 1.315 4.94 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2525 0.7025 0.4375 0.7025 0.4375 0.2125 0.5025 0.2125 0.5025 1.2375 0.4375 1.2375 0.4375 0.8375 0.2525 0.8375  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.9525 0.5425 4.57 0.5425 4.57 0.6075 4.1175 0.6075 4.1175 0.6975 4.0525 0.6975 4.0525 0.6425 3.9525 0.6425  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 4.94 -0.085 4.94 0.085 4.64 0.085 4.64 0.1925 4.575 0.1925 4.575 0.085 3.8225 0.085 3.8225 0.1925 3.7575 0.1925 3.7575 0.085 3.4775 0.085 3.4775 0.1925 3.4125 0.1925 3.4125 0.085 2.7525 0.085 2.7525 0.235 2.6175 0.235 2.6175 0.085 1.8825 0.085 1.8825 0.1925 1.8175 0.1925 1.8175 0.085 0.9175 0.085 0.9175 0.27 0.8525 0.27 0.8525 0.085 0.3125 0.085 0.3125 0.2425 0.2475 0.2425 0.2475 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.8625 0.7025 3.9275 0.7025 3.9275 0.8425 4.4125 0.8425 4.4125 0.9225 4.5925 0.9225 4.5925 0.9875 4.3475 0.9875 4.3475 0.9075 3.8625 0.9075  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.4825 0.7025 3.5475 0.7025 3.5475 0.8375 3.4825 0.8375  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.5725 0.3725 0.6475 0.3725 0.6475 0.1625 0.7125 0.1625 0.7125 0.4375 0.6375 0.4375 0.6375 1.115 0.6575 1.115 0.6575 1.25 0.5725 1.25  ;
        POLYGON 1.17 1.1125 1.9825 1.1125 1.9825 1.2475 1.9175 1.2475 1.9175 1.1775 1.2225 1.1775 1.2225 1.25 1.1575 1.25 1.1575 1.1775 1.105 1.1775 1.105 0.5275 0.8375 0.5275 0.8375 0.8025 0.7025 0.8025 0.7025 0.7375 0.7725 0.7375 0.7725 0.4625 1.105 0.4625 1.105 0.22 1.4175 0.22 1.4175 0.15 1.4825 0.15 1.4825 0.285 1.17 0.285  ;
        POLYGON 2.2775 0.15 2.3425 0.15 2.3425 0.31 2.8125 0.31 2.8125 0.375 2.2775 0.375  ;
        POLYGON 2.4525 0.9925 2.4775 0.9925 2.4775 0.98 2.8125 0.98 2.8125 1.045 2.5175 1.045 2.5175 1.25 2.4525 1.25  ;
        POLYGON 1.235 0.35 2.0025 0.35 2.0025 0.1625 2.0675 0.1625 2.0675 0.44 2.9675 0.44 2.9675 0.505 2.0025 0.505 2.0025 0.415 1.3 0.415 1.3 0.9825 2.1375 0.9825 2.1375 1.2375 2.0725 1.2375 2.0725 1.0475 1.235 1.0475  ;
        POLYGON 1.7125 0.5725 3.0325 0.5725 3.0325 0.15 3.0975 0.15 3.0975 0.6125 3.1025 0.6125 3.1025 1.12 3.0375 1.12 3.0375 0.6375 1.7125 0.6375  ;
        POLYGON 3.2325 0.96 3.6675 0.96 3.6675 1.12 3.6025 1.12 3.6025 1.025 3.2325 1.025 3.2325 1.25 2.9075 1.25 2.9075 0.92 2.8375 0.92 2.8375 0.785 1.5825 0.785 1.5825 0.545 1.365 0.545 1.365 0.48 1.6475 0.48 1.6475 0.72 2.9025 0.72 2.9025 0.855 2.9725 0.855 2.9725 1.185 3.1675 1.185 3.1675 0.2575 3.6025 0.2575 3.6025 0.1625 3.6675 0.1625 3.6675 0.3225 3.2325 0.3225  ;
        POLYGON 3.7975 0.9725 4.2825 0.9725 4.2825 1.1475 4.2175 1.1475 4.2175 1.0375 3.7325 1.0375 3.7325 0.6375 3.2975 0.6375 3.2975 0.5725 3.7325 0.5725 3.7325 0.3225 3.7375 0.3225 3.7375 0.2825 4.1925 0.2825 4.1925 0.1625 4.2575 0.1625 4.2575 0.3475 3.7975 0.3475  ;
        POLYGON 4.0775 0.4125 4.765 0.4125 4.765 0.1625 4.83 0.1625 4.83 0.4275 4.8525 0.4275 4.8525 1.1475 4.7875 1.1475 4.7875 0.4775 4.0775 0.4775  ;
  END
END SDFFR_X2

MACRO SDFFS_X1
  CLASS core ;
  FOREIGN SDFFS_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 5.13 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 4.5775 0.3775 4.6425 0.3775 4.6425 0.5625 4.6875 0.5625 4.6875 0.6975 4.6425 0.6975 4.6425 0.8375 4.5775 0.8375  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.92 0.3475 3.8025 0.3475 3.8025 0.365 4.1175 0.365 4.1175 0.5575 4.0525 0.5575 4.0525 0.43 3.7575 0.43 3.7575 0.4125 2.985 0.4125 2.985 0.4825 2.92 0.4825  ;
    END
  END SN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1925 0.3875 0.2575 0.3875 0.2575 0.4575 0.3525 0.4575 0.3525 0.5225 0.1925 0.5225 0.1925 0.4575  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2475 1.315 0.2475 0.9775 0.3125 0.9775 0.3125 1.315 1.0075 1.315 1.0075 0.9775 1.0725 0.9775 1.0725 1.315 1.5125 1.315 1.5125 0.9725 1.5775 0.9725 1.5775 1.315 1.8425 1.315 1.8425 1.2 1.9075 1.2 1.9075 1.315 2.6175 1.315 2.6175 1.1125 2.6825 1.1125 2.6825 1.315 3.23 1.315 3.23 1.1075 3.295 1.1075 3.295 1.315 4.05 1.315 4.05 0.9525 4.115 0.9525 4.115 1.315 4.425 1.315 4.425 0.9125 4.49 0.9125 4.49 1.315 4.7625 1.315 4.7625 0.7625 4.8275 0.7625 4.8275 1.315 5.13 1.315 5.13 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 4.8125 0.5625 4.9525 0.5625 4.9525 0.3775 5.0175 0.3775 5.0175 0.8375 4.9525 0.8375 4.9525 0.6975 4.8125 0.6975  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3625 0.3225 0.4425 0.3225 0.4425 0.2825 0.5325 0.2825 0.5325 0.3875 0.9275 0.3875 0.9275 0.5225 0.8625 0.5225 0.8625 0.4525 0.4425 0.4525 0.4425 0.3875 0.3625 0.3875  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 5.13 -0.085 5.13 0.085 4.8275 0.085 4.8275 0.4975 4.7625 0.4975 4.7625 0.085 4.1275 0.085 4.1275 0.3 3.9925 0.3 3.9925 0.085 3.125 0.085 3.125 0.2825 2.99 0.2825 2.99 0.085 2.0325 0.085 2.0325 0.3175 1.9675 0.3175 1.9675 0.085 1.6175 0.085 1.6175 0.1925 1.5525 0.1925 1.5525 0.085 1.1575 0.085 1.1575 0.1925 1.0925 0.1925 1.0925 0.085 0.3125 0.085 0.3125 0.1925 0.2475 0.1925 0.2475 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3225 0.7175 0.9875 0.7175 0.9875 0.6475 1.0525 0.6475 1.0525 0.7825 0.5075 0.7825 0.5075 0.9775 0.4425 0.9775 0.4425 0.7825 0.3225 0.7825  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.3575 0.4575 1.4475 0.4575 1.5125 0.4575 1.5125 0.48 1.5475 0.48 1.5475 0.545 1.5125 0.545 1.51 0.545 1.4475 0.545 1.3575 0.545  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.0625 0.1625 0.1275 0.1625 0.1275 0.5875 0.7125 0.5875 0.7125 0.5175 0.7775 0.5175 0.7775 0.6525 0.1275 0.6525 0.1275 1.0575 0.0625 1.0575  ;
        POLYGON 1.2475 0.7775 1.3825 0.7775 1.3825 0.925 1.4275 0.925 1.4275 0.99 1.2925 0.99 1.2925 0.8425 1.2475 0.8425  ;
        POLYGON 1.4325 0.3225 1.5975 0.3225 1.5975 0.2875 1.6625 0.2875 1.6625 0.4225 1.5975 0.4225 1.5975 0.3875 1.3675 0.3875 1.2725 0.3875 1.2725 0.3225 1.3675 0.3225 1.3675 0.215 1.3325 0.215 1.3325 0.15 1.4675 0.15 1.4675 0.215 1.4325 0.215  ;
        POLYGON 1.7425 0.1625 1.8125 0.1625 1.8125 0.5475 1.7425 0.5475  ;
        POLYGON 1.7025 0.7625 1.8475 0.7625 1.8475 0.8275 1.7675 0.8275 1.7675 1.0025 1.7025 1.0025  ;
        POLYGON 0.5975 0.9575 0.6675 0.9575 0.6675 0.8475 1.1175 0.8475 1.1175 0.3225 0.6975 0.3225 0.6975 0.3125 0.6675 0.3125 0.6675 0.2625 0.5975 0.2625 0.5975 0.1975 0.7325 0.1975 0.7325 0.2575 1.1825 0.2575 1.1825 0.6125 1.9225 0.6125 1.9225 0.4625 1.9875 0.4625 1.9875 0.8725 1.9225 0.8725 1.9225 0.6775 1.1825 0.6775 1.1825 0.9125 0.7325 0.9125 0.7325 1.0225 0.5975 1.0225  ;
        POLYGON 2.2425 0.4625 2.3075 0.4625 2.3075 0.7375 2.9875 0.7375 2.9875 0.8025 2.3675 0.8025 2.3675 0.8725 2.26 0.8725 2.26 0.7825 2.2425 0.7825  ;
        POLYGON 2.5725 0.5375 2.6375 0.5375 2.6375 0.5475 3.12 0.5475 3.12 0.4775 3.185 0.4775 3.185 0.5475 3.2325 0.5475 3.2325 0.9125 3.1675 0.9125 3.1675 0.6125 2.6375 0.6125 2.6375 0.6725 2.5725 0.6725  ;
        POLYGON 2.1775 0.9825 2.9925 0.9825 2.9925 0.9125 3.0575 0.9125 3.0575 0.9775 3.2975 0.9775 3.2975 0.5275 3.3725 0.5275 3.3725 1.0125 3.3525 1.0125 3.3525 1.0425 3.0575 1.0425 3.0575 1.0475 2.3175 1.0475 2.3175 1.195 2.1825 1.195 2.1825 1.0475 2.1175 1.0475 2.1175 1.0075 2.1125 1.0075 2.1125 0.2675 2.3425 0.2675 2.3425 0.1975 2.4075 0.1975 2.4075 0.3325 2.1775 0.3325  ;
        POLYGON 3.4475 0.4775 3.5125 0.4775 3.5125 0.7875 3.73 0.7875 3.73 0.8525 3.4475 0.8525  ;
        POLYGON 3.62 1.0375 3.79 1.0375 3.79 0.8775 3.795 0.8775 3.795 0.6475 3.6475 0.6475 3.6475 0.5425 3.5775 0.5425 3.5775 0.4775 3.7125 0.4775 3.7125 0.5825 3.855 0.5825 3.855 0.6225 4.38 0.6225 4.38 0.6875 3.86 0.6875 3.86 0.9025 3.855 0.9025 3.855 1.1025 3.62 1.1025  ;
        POLYGON 4.005 0.7525 4.445 0.7525 4.445 0.535 4.4375 0.535 4.4375 0.355 4.3675 0.355 4.3675 0.15 4.5025 0.15 4.5025 0.5025 4.5125 0.5025 4.5125 0.6375 4.51 0.6375 4.51 0.8175 4.3 0.8175 4.3 1.0325 4.235 1.0325 4.235 0.8875 4.005 0.8875  ;
  END
END SDFFS_X1

MACRO SDFFS_X2
  CLASS core ;
  FOREIGN SDFFS_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 5.13 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 4.5775 0.3775 4.665 0.3775 4.665 0.5625 4.6875 0.5625 4.6875 0.6975 4.665 0.6975 4.665 0.8375 4.5775 0.8375  ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.92 0.3475 3.8025 0.3475 3.8025 0.365 4.1175 0.365 4.1175 0.5575 4.0525 0.5575 4.0525 0.43 3.7575 0.43 3.7575 0.4125 2.985 0.4125 2.985 0.4825 2.92 0.4825  ;
    END
  END SN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1925 0.3875 0.2575 0.3875 0.2575 0.4575 0.3525 0.4575 0.3525 0.5225 0.1925 0.5225 0.1925 0.4575  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2475 1.315 0.2475 0.9775 0.3125 0.9775 0.3125 1.315 1.0075 1.315 1.0075 0.9775 1.0725 0.9775 1.0725 1.315 1.5125 1.315 1.5125 0.9725 1.5775 0.9725 1.5775 1.315 1.8425 1.315 1.8425 1.2 1.9075 1.2 1.9075 1.315 2.6175 1.315 2.6175 1.1125 2.6825 1.1125 2.6825 1.315 3.23 1.315 3.23 1.1075 3.295 1.1075 3.295 1.315 4.05 1.315 4.05 0.9525 4.115 0.9525 4.115 1.315 4.425 1.315 4.425 0.9125 4.49 0.9125 4.49 1.315 4.785 1.315 4.785 0.7625 4.85 0.7625 4.85 1.315 5.13 1.315 5.13 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 4.8125 0.5625 4.9525 0.5625 4.9525 0.3775 5.04 0.3775 5.04 0.8375 4.9525 0.8375 4.9525 0.6975 4.8125 0.6975  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3625 0.3225 0.4425 0.3225 0.4425 0.2825 0.5325 0.2825 0.5325 0.3875 0.9275 0.3875 0.9275 0.5225 0.8625 0.5225 0.8625 0.4525 0.4425 0.4525 0.4425 0.3875 0.3625 0.3875  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 5.13 -0.085 5.13 0.085 4.85 0.085 4.85 0.4975 4.785 0.4975 4.785 0.085 4.1275 0.085 4.1275 0.3 3.9925 0.3 3.9925 0.085 3.125 0.085 3.125 0.2825 2.99 0.2825 2.99 0.085 2.0325 0.085 2.0325 0.3175 1.9675 0.3175 1.9675 0.085 1.6175 0.085 1.6175 0.1925 1.5525 0.1925 1.5525 0.085 1.1575 0.085 1.1575 0.1925 1.0925 0.1925 1.0925 0.085 0.3125 0.085 0.3125 0.1925 0.2475 0.1925 0.2475 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3225 0.7175 0.9875 0.7175 0.9875 0.6475 1.0525 0.6475 1.0525 0.7825 0.5075 0.7825 0.5075 0.9775 0.4425 0.9775 0.4425 0.7825 0.3225 0.7825  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.3575 0.4575 1.4475 0.4575 1.5125 0.4575 1.5125 0.48 1.5475 0.48 1.5475 0.545 1.5125 0.545 1.51 0.545 1.4475 0.545 1.3575 0.545  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.0625 0.1625 0.1275 0.1625 0.1275 0.5875 0.7125 0.5875 0.7125 0.5175 0.7775 0.5175 0.7775 0.6525 0.1275 0.6525 0.1275 1.0575 0.0625 1.0575  ;
        POLYGON 1.2475 0.7775 1.3825 0.7775 1.3825 0.925 1.4275 0.925 1.4275 0.99 1.2925 0.99 1.2925 0.8425 1.2475 0.8425  ;
        POLYGON 1.4325 0.3225 1.5975 0.3225 1.5975 0.2875 1.6625 0.2875 1.6625 0.4225 1.5975 0.4225 1.5975 0.3875 1.3675 0.3875 1.2725 0.3875 1.2725 0.3225 1.3675 0.3225 1.3675 0.215 1.3325 0.215 1.3325 0.15 1.4675 0.15 1.4675 0.215 1.4325 0.215  ;
        POLYGON 1.7425 0.1625 1.8125 0.1625 1.8125 0.5475 1.7425 0.5475  ;
        POLYGON 1.7025 0.7625 1.8475 0.7625 1.8475 0.8275 1.7675 0.8275 1.7675 1.0025 1.7025 1.0025  ;
        POLYGON 0.5975 0.9575 0.6675 0.9575 0.6675 0.8475 1.1175 0.8475 1.1175 0.3225 0.6975 0.3225 0.6975 0.3125 0.6675 0.3125 0.6675 0.2625 0.5975 0.2625 0.5975 0.1975 0.7325 0.1975 0.7325 0.2575 1.1825 0.2575 1.1825 0.6125 1.9225 0.6125 1.9225 0.4625 1.9875 0.4625 1.9875 0.8725 1.9225 0.8725 1.9225 0.6775 1.1825 0.6775 1.1825 0.9125 0.7325 0.9125 0.7325 1.0225 0.5975 1.0225  ;
        POLYGON 2.2425 0.4625 2.3075 0.4625 2.3075 0.7375 2.9875 0.7375 2.9875 0.8025 2.3675 0.8025 2.3675 0.8725 2.26 0.8725 2.26 0.7825 2.2425 0.7825  ;
        POLYGON 2.5725 0.5375 2.6375 0.5375 2.6375 0.5475 3.12 0.5475 3.12 0.4775 3.185 0.4775 3.185 0.5475 3.2325 0.5475 3.2325 0.9125 3.1675 0.9125 3.1675 0.6125 2.6375 0.6125 2.6375 0.6725 2.5725 0.6725  ;
        POLYGON 2.1775 0.9825 2.9925 0.9825 2.9925 0.9125 3.0575 0.9125 3.0575 0.9775 3.2975 0.9775 3.2975 0.5275 3.3725 0.5275 3.3725 1.0125 3.3525 1.0125 3.3525 1.0425 3.0575 1.0425 3.0575 1.0475 2.3175 1.0475 2.3175 1.195 2.1825 1.195 2.1825 1.0475 2.1175 1.0475 2.1175 1.0075 2.1125 1.0075 2.1125 0.2675 2.3425 0.2675 2.3425 0.1975 2.4075 0.1975 2.4075 0.3325 2.1775 0.3325  ;
        POLYGON 3.4475 0.4775 3.5125 0.4775 3.5125 0.7875 3.73 0.7875 3.73 0.8525 3.4475 0.8525  ;
        POLYGON 3.62 1.0375 3.79 1.0375 3.79 0.8775 3.795 0.8775 3.795 0.6475 3.6475 0.6475 3.6475 0.5425 3.5775 0.5425 3.5775 0.4775 3.7125 0.4775 3.7125 0.5825 3.855 0.5825 3.855 0.6225 4.38 0.6225 4.38 0.6875 3.86 0.6875 3.86 0.9025 3.855 0.9025 3.855 1.1025 3.62 1.1025  ;
        POLYGON 4.005 0.7525 4.445 0.7525 4.445 0.355 4.3675 0.355 4.3675 0.15 4.5125 0.15 4.5125 0.6375 4.51 0.6375 4.51 0.8175 4.3 0.8175 4.3 1.0325 4.235 1.0325 4.235 0.8875 4.005 0.8875  ;
  END
END SDFFS_X2

MACRO SDFF_X1
  CLASS core ;
  FOREIGN SDFF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 4.37 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4375 0.1975 0.5075 0.1975 0.5075 1.25 0.4375 1.25  ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.7575 0.7125 3.9975 0.7125 3.9975 0.7375 4.1525 0.7375 4.1525 0.8025 3.9325 0.8025 3.9325 0.7775 3.7575 0.7775  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2475 1.315 0.2475 1.17 0.3125 1.17 0.3125 1.315 0.7775 1.315 0.7775 1.13 0.8425 1.13 0.8425 1.315 1.5375 1.315 1.5375 1.2075 1.6025 1.2075 1.6025 1.315 2.1025 1.315 2.1025 1.18 2.1675 1.18 2.1675 1.315 2.8825 1.315 2.8825 1.18 2.9475 1.18 2.9475 1.185 3.3075 1.185 3.3075 1.17 3.3725 1.17 3.3725 1.185 4.0625 1.185 4.0625 1.03 4.1275 1.03 4.1275 1.315 4.37 1.315 4.37 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.1975 0.1275 0.1975 0.1275 1.25 0.0625 1.25  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.4175 0.5625 4.035 0.5625 4.035 0.6275 3.5525 0.6275 3.5525 0.6975 3.4825 0.6975 3.4825 0.665 3.4175 0.665  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 4.37 -0.085 4.37 0.085 4.105 0.085 4.105 0.1925 4.04 0.1925 4.04 0.085 3.2875 0.085 3.2875 0.1925 3.2225 0.1925 3.2225 0.085 2.9225 0.085 2.9225 0.1925 2.8575 0.1925 2.8575 0.085 2.1625 0.085 2.1625 0.27 2.0975 0.27 2.0975 0.085 1.6025 0.085 1.6025 0.3175 1.5375 0.3175 1.5375 0.085 0.8425 0.085 0.8425 0.3175 0.7775 0.3175 0.7775 0.085 0.3125 0.085 0.3125 0.3175 0.2475 0.3175 0.2475 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.3275 0.725 3.3925 0.725 3.3925 0.8425 3.8775 0.8425 3.8775 0.8775 4.0575 0.8775 4.0575 0.95 3.8125 0.95 3.8125 0.9075 3.3275 0.9075  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.9125 0.7025 2.9775 0.7025 2.9775 0.7725 3.0625 0.7725 3.0625 0.8375 2.9125 0.8375  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.5925 0.1625 0.6575 0.1625 0.6575 1.25 0.5925 1.25  ;
        POLYGON 0.7875 1 0.9725 1 0.9725 1.115 1.2225 1.115 1.2225 1.25 1.1575 1.25 1.1575 1.18 0.9075 1.18 0.9075 1.065 0.7225 1.065 0.7225 0.415 0.7525 0.415 0.7525 0.405 1.1575 0.405 1.1575 0.1975 1.2225 0.1975 1.2225 0.47 0.7875 0.47  ;
        POLYGON 1.8675 0.2225 1.9125 0.2225 1.9125 0.15 1.9775 0.15 1.9775 0.285 1.9325 0.285 1.9325 0.425 1.8675 0.425  ;
        POLYGON 1.8575 0.87 2.2875 0.87 2.2875 0.935 1.9475 0.935 1.9475 1.25 1.8825 1.25 1.8825 0.935 1.8575 0.935  ;
        POLYGON 1.0375 0.985 1.1425 0.985 1.1425 0.535 1.7275 0.535 1.7275 0.2875 1.7925 0.2875 1.7925 0.535 2.4725 0.535 2.4725 0.6 1.2075 0.6 1.2075 0.985 1.3175 0.985 1.3175 1.005 1.7925 1.005 1.7925 1.2375 1.7275 1.2375 1.7275 1.07 1.27 1.07 1.27 1.05 1.0375 1.05  ;
        POLYGON 2.04 0.335 2.2275 0.335 2.2275 0.22 2.4775 0.22 2.4775 0.15 2.5425 0.15 2.5425 0.285 2.2925 0.285 2.2925 0.4 2.105 0.4 2.105 0.47 2.04 0.47  ;
        POLYGON 2.0125 1.05 2.2725 1.05 2.2725 1.075 2.5675 1.075 2.5675 1.21 2.5025 1.21 2.5025 1.14 2.22 1.14 2.22 1.115 2.0125 1.115  ;
        POLYGON 2.6175 0.945 3.1325 0.945 3.1325 1.12 3.0675 1.12 3.0675 1.01 2.3675 1.01 2.3675 0.945 2.5525 0.945 2.5525 0.75 1.2725 0.75 1.2725 0.685 2.5525 0.685 2.5525 0.35 2.6225 0.35 2.6225 0.2575 3.0475 0.2575 3.0475 0.1625 3.1125 0.1625 3.1125 0.3225 2.6875 0.3225 2.6875 0.415 2.6175 0.415  ;
        POLYGON 3.2625 0.975 3.7475 0.975 3.7475 1.11 3.6825 1.11 3.6825 1.04 3.1975 1.04 3.1975 0.6375 2.7425 0.6375 2.7425 0.5725 3.1975 0.5725 3.1975 0.3275 3.21 0.3275 3.21 0.3025 3.635 0.3025 3.635 0.1625 3.7 0.1625 3.7 0.3675 3.2625 0.3675  ;
        POLYGON 3.5425 0.4325 4.23 0.4325 4.23 0.1625 4.295 0.1625 4.295 0.4475 4.3175 0.4475 4.3175 1.25 4.2525 1.25 4.2525 0.4975 3.5425 0.4975  ;
  END
END SDFF_X1

MACRO SDFF_X2
  CLASS core ;
  FOREIGN SDFF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 4.37 BY 1.4 ;
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4375 0.1975 0.5075 0.1975 0.5075 1.25 0.4375 1.25  ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.7575 0.7125 3.9975 0.7125 3.9975 0.7375 4.1525 0.7375 4.1525 0.8025 3.9325 0.8025 3.9325 0.7775 3.7575 0.7775  ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2475 1.315 0.2475 1.03 0.3125 1.03 0.3125 1.315 0.7775 1.315 0.7775 1.13 0.8425 1.13 0.8425 1.315 1.5375 1.315 1.5375 1.2075 1.6025 1.2075 1.6025 1.315 2.1025 1.315 2.1025 1.18 2.1675 1.18 2.1675 1.315 2.8825 1.315 2.8825 1.18 2.9475 1.18 2.9475 1.185 3.3075 1.185 3.3075 1.17 3.3725 1.17 3.3725 1.185 4.0625 1.185 4.0625 1.03 4.1275 1.03 4.1275 1.315 4.37 1.315 4.37 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.0625 0.2125 0.1275 0.2125 0.1275 1.11 0.0625 1.11  ;
    END
  END Q
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.4175 0.5625 4.035 0.5625 4.035 0.6275 3.5525 0.6275 3.5525 0.6975 3.4825 0.6975 3.4825 0.665 3.4175 0.665  ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 4.37 -0.085 4.37 0.085 4.105 0.085 4.105 0.1925 4.04 0.1925 4.04 0.085 3.2875 0.085 3.2875 0.1925 3.2225 0.1925 3.2225 0.085 2.9225 0.085 2.9225 0.1925 2.8575 0.1925 2.8575 0.085 2.1625 0.085 2.1625 0.27 2.0975 0.27 2.0975 0.085 1.6025 0.085 1.6025 0.3175 1.5375 0.3175 1.5375 0.085 0.8425 0.085 0.8425 0.3175 0.7775 0.3175 0.7775 0.085 0.3125 0.085 0.3125 0.3175 0.2475 0.3175 0.2475 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 3.3275 0.725 3.3925 0.725 3.3925 0.8425 3.8775 0.8425 3.8775 0.8775 4.0575 0.8775 4.0575 0.9425 3.8125 0.9425 3.8125 0.9075 3.3275 0.9075  ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.9125 0.7025 2.9775 0.7025 2.9775 0.7725 3.0625 0.7725 3.0625 0.8375 2.9125 0.8375  ;
    END
  END CK
  OBS
      LAYER metal1 ;
        POLYGON 0.5925 0.1625 0.6575 0.1625 0.6575 1.25 0.5925 1.25  ;
        POLYGON 0.7875 1 0.9725 1 0.9725 1.115 1.2225 1.115 1.2225 1.25 1.1575 1.25 1.1575 1.18 0.9075 1.18 0.9075 1.065 0.7225 1.065 0.7225 0.415 0.7525 0.415 0.7525 0.405 1.1575 0.405 1.1575 0.1975 1.2225 0.1975 1.2225 0.47 0.7875 0.47  ;
        POLYGON 1.8675 0.2225 1.9125 0.2225 1.9125 0.15 1.9775 0.15 1.9775 0.285 1.9325 0.285 1.9325 0.425 1.8675 0.425  ;
        POLYGON 1.8575 0.87 2.2875 0.87 2.2875 0.935 1.9475 0.935 1.9475 1.25 1.8825 1.25 1.8825 0.935 1.8575 0.935  ;
        POLYGON 1.0375 0.985 1.1425 0.985 1.1425 0.535 1.7275 0.535 1.7275 0.2875 1.7925 0.2875 1.7925 0.535 2.4725 0.535 2.4725 0.6 1.2075 0.6 1.2075 0.985 1.3175 0.985 1.3175 1.005 1.7925 1.005 1.7925 1.2375 1.7275 1.2375 1.7275 1.07 1.27 1.07 1.27 1.05 1.0375 1.05  ;
        POLYGON 2.04 0.335 2.2275 0.335 2.2275 0.22 2.4775 0.22 2.4775 0.15 2.5425 0.15 2.5425 0.285 2.2925 0.285 2.2925 0.4 2.105 0.4 2.105 0.47 2.04 0.47  ;
        POLYGON 2.0125 1.05 2.2725 1.05 2.2725 1.075 2.5675 1.075 2.5675 1.21 2.5025 1.21 2.5025 1.14 2.22 1.14 2.22 1.115 2.0125 1.115  ;
        POLYGON 2.6175 0.945 3.1325 0.945 3.1325 1.12 3.0675 1.12 3.0675 1.01 2.3675 1.01 2.3675 0.945 2.5525 0.945 2.5525 0.75 1.2725 0.75 1.2725 0.685 2.5525 0.685 2.5525 0.35 2.6225 0.35 2.6225 0.2575 3.0475 0.2575 3.0475 0.1625 3.1125 0.1625 3.1125 0.3225 2.6875 0.3225 2.6875 0.415 2.6175 0.415  ;
        POLYGON 3.2625 0.975 3.7475 0.975 3.7475 1.11 3.6825 1.11 3.6825 1.04 3.1975 1.04 3.1975 0.6375 2.7425 0.6375 2.7425 0.5725 3.1975 0.5725 3.1975 0.3275 3.21 0.3275 3.21 0.3025 3.635 0.3025 3.635 0.1625 3.7 0.1625 3.7 0.3675 3.2625 0.3675  ;
        POLYGON 3.5425 0.4325 4.23 0.4325 4.23 0.1625 4.295 0.1625 4.295 0.4475 4.3175 0.4475 4.3175 1.25 4.2525 1.25 4.2525 0.4975 3.5425 0.4975  ;
  END
END SDFF_X2

MACRO TBUF_X1
  CLASS core ;
  FOREIGN TBUF_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.5625 0.6375 0.5625 0.6375 0.2725 0.7025 0.2725 0.7025 0.79 0.6375 0.79 0.6375 0.6975 0.6325 0.6975  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1825 0.565 0.2525 0.565 0.2525 0.5625 0.3175 0.5625 0.3175 0.6975 0.1825 0.6975  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2075 1.315 0.2075 0.815 0.3425 0.815 0.3425 1.315 0.9875 1.315 0.9875 0.9725 1.0525 0.9725 1.0525 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 1.0625 0.085 1.0625 0.35 0.9975 0.35 0.9975 0.085 0.3625 0.085 0.3625 0.3175 0.2275 0.3175 0.2275 0.085 0 0.085  ;
    END
  END VSS
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.0125 0.5625 1.0775 0.5625 1.0775 0.6975 1.0125 0.6975  ;
    END
  END EN
  OBS
      LAYER metal1 ;
        POLYGON 0.7675 0.27 0.9125 0.27 0.9125 0.335 0.8325 0.335 0.8325 0.9475 0.9025 0.9475 0.9025 1.0125 0.7675 1.0125  ;
        POLYGON 0.0525 0.4725 0.0575 0.4725 0.0575 0.2725 0.1225 0.2725 0.1225 0.4325 0.4425 0.4325 0.4425 0.4975 0.1175 0.4975 0.1175 0.855 0.0525 0.855  ;
  END
END TBUF_X1

MACRO TBUF_X16
  CLASS core ;
  FOREIGN TBUF_X16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 3.61 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.695 0.94 0.74 0.94 0.74 1.08 1.43 1.08 1.43 1.005 1.365 1.005 1.365 0.94 2.255 0.94 2.255 1.08 2.8775 1.08 2.8775 0.94 3.015 0.94 3.015 1.145 2.125 1.145 2.125 1.08 2.19 1.08 2.19 1.005 1.495 1.005 1.495 1.145 0.605 1.145 0.605 0.94 0.63 0.94 0.63 0.3675 0.605 0.3675 0.605 0.1625 0.74 0.1625 0.74 0.3875 1.36 0.3875 1.36 0.1625 1.495 0.1625 1.495 0.3875 2.12 0.3875 2.12 0.1625 2.255 0.1625 2.255 0.3875 2.88 0.3875 2.88 0.1625 3.015 0.1625 3.015 0.3675 2.945 0.3675 2.945 0.4525 0.695 0.4525  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.185 0.5275 0.25 0.5275 0.25 0.5975 0.3525 0.5975 0.3525 0.6625 0.185 0.6625  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.26 1.315 0.26 1.0675 0.325 1.0675 0.325 1.315 0.98 1.315 0.98 1.2425 1.115 1.2425 1.115 1.315 1.74 1.315 1.74 1.1025 1.875 1.1025 1.875 1.315 2.5 1.315 2.5 1.2425 2.635 1.2425 2.635 1.315 3.295 1.315 3.295 1.0675 3.36 1.0675 3.36 1.315 3.61 1.315 3.61 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 3.61 -0.085 3.61 0.085 3.36 0.085 3.36 0.3575 3.295 0.3575 3.295 0.085 2.635 0.085 2.635 0.3225 2.5 0.3225 2.5 0.085 1.875 0.085 1.875 0.3225 1.74 0.3225 1.74 0.085 1.115 0.085 1.115 0.3225 0.98 0.3225 0.98 0.085 0.36 0.085 0.36 0.3225 0.225 0.3225 0.225 0.085 0 0.085  ;
    END
  END VSS
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.785 0.6675 3.37 0.6675 3.37 0.5975 3.435 0.5975 3.435 0.7325 0.9225 0.7325 0.9225 0.8025 0.85 0.8025 0.85 0.8925 0.785 0.8925  ;
    END
  END EN
  OBS
      LAYER metal1 ;
        POLYGON 1.09 0.7975 3.29 0.7975 3.29 0.8625 1.09 0.8625  ;
        POLYGON 0.76 0.5175 3.025 0.5175 3.025 0.4475 3.5 0.4475 3.5 0.2675 3.565 0.2675 3.565 1.0225 3.5 1.0225 3.5 0.5125 3.09 0.5125 3.09 0.5825 0.76 0.5825  ;
        POLYGON 0.055 0.2675 0.12 0.2675 0.12 0.7625 0.405 0.7625 0.405 0.8975 0.34 0.8975 0.34 0.8275 0.12 0.8275 0.12 1.0225 0.055 1.0225  ;
  END
END TBUF_X16

MACRO TBUF_X2
  CLASS core ;
  FOREIGN TBUF_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.2075 0.6975 0.2075 0.6975 1.1025 0.6325 1.1025  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2125 0.7025 0.3175 0.7025 0.3175 0.8375 0.2125 0.8375  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2575 1.315 0.2575 1.0075 0.3225 1.0075 0.3225 1.315 0.9725 1.315 0.9725 0.8525 1.0375 0.8525 1.0375 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 1.0375 0.085 1.0375 0.3575 0.9725 0.3575 0.9725 0.085 0.3225 0.085 0.3225 0.4375 0.2575 0.4375 0.2575 0.085 0 0.085  ;
    END
  END VSS
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.0125 0.4225 1.0775 0.4225 1.0775 0.5575 1.0125 0.5575  ;
    END
  END EN
  OBS
      LAYER metal1 ;
        POLYGON 0.7875 0.2425 0.8525 0.2425 0.8525 0.9275 0.7875 0.9275  ;
        POLYGON 0.0525 0.3475 0.1175 0.3475 0.1175 0.5725 0.3375 0.5725 0.3375 0.5025 0.4025 0.5025 0.4025 0.6375 0.1175 0.6375 0.1175 1.2225 0.0525 1.2225  ;
  END
END TBUF_X2

MACRO TBUF_X4
  CLASS core ;
  FOREIGN TBUF_X4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.33 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.5975 0.1725 0.7375 0.1725 0.7375 0.2375 0.6975 0.2375 0.6975 0.2775 0.6975 0.3975 0.6975 1.12 0.6325 1.12 0.6325 0.3975 0.6325 0.2775 0.6325 0.2375 0.5975 0.2375  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2075 0.7025 0.3175 0.7025 0.3175 0.8375 0.2075 0.8375  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2525 1.315 0.2525 1.025 0.3175 1.025 0.3175 1.315 1.0075 1.315 1.0075 1.0675 1.0725 1.0675 1.0725 1.315 1.33 1.315 1.33 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.33 -0.085 1.33 0.085 1.0725 0.085 1.0725 0.3675 1.0075 0.3675 1.0075 0.085 0.3175 0.085 0.3175 0.38 0.2525 0.38 0.2525 0.085 0 0.085  ;
    END
  END VSS
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.7775 0.6325 1.0125 0.6325 1.0125 0.5625 1.1175 0.5625 1.1175 0.6975 0.8425 0.6975 0.8425 0.7675 0.7775 0.7675  ;
    END
  END EN
  OBS
      LAYER metal1 ;
        POLYGON 0.7775 0.4325 1.2125 0.4325 1.2125 0.2775 1.2775 0.2775 1.2775 1.0225 1.2125 1.0225 1.2125 0.4975 0.8425 0.4975 0.8425 0.5675 0.7775 0.5675  ;
        POLYGON 0.0475 0.2775 0.1125 0.2775 0.1125 0.385 0.1125 0.39 0.1125 0.57 0.4475 0.57 0.4475 0.635 0.4475 1.185 0.8775 1.185 0.8775 0.8425 0.9075 0.8425 0.9075 0.7625 0.9725 0.7625 0.9725 0.8975 0.9425 0.8975 0.9425 1.25 0.3825 1.25 0.3825 0.635 0.1125 0.635 0.1125 1.24 0.0475 1.24 0.0475 0.635 0.0475 0.57 0.0475 0.39 0.0475 0.385  ;
  END
END TBUF_X4

MACRO TBUF_X8
  CLASS core ;
  FOREIGN TBUF_X8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.28 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.4975 1.0225 1.5275 1.0225 1.5275 1.0875 1.3925 1.0875 1.3925 1.0225 1.4325 1.0225 1.4325 0.4525 0.7025 0.4525 0.7025 1.03 0.7375 1.03 0.7375 1.095 0.6025 1.095 0.6025 1.03 0.6375 1.03 0.6375 0.3675 0.6225 0.3675 0.6225 0.1625 0.7575 0.1625 0.7575 0.3875 1.3575 0.3875 1.3575 0.3175 1.3775 0.3175 1.3775 0.1625 1.5125 0.1625 1.5125 0.3675 1.4975 0.3675  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1825 0.765 0.3175 0.765 0.3175 0.9775 0.2525 0.9775 0.2525 0.83 0.1825 0.83  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.2275 1.315 0.2275 1.07 0.3625 1.07 0.3625 1.315 0.9975 1.315 0.9975 1.2425 1.1325 1.2425 1.1325 1.315 1.7725 1.315 1.7725 1.0625 1.9075 1.0625 1.9075 1.315 2.28 1.315 2.28 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.28 -0.085 2.28 0.085 1.9275 0.085 1.9275 0.3225 1.7925 0.3225 1.7925 0.085 1.1325 0.085 1.1325 0.3225 0.9975 0.3225 0.9975 0.085 0.3775 0.085 0.3775 0.3225 0.2425 0.3225 0.2425 0.085 0 0.085  ;
    END
  END VSS
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.7675 0.6675 1.3675 0.6675 1.3675 0.7325 1.3025 0.7325 1.3025 0.8025 1.1675 0.8025 1.1675 0.7325 0.7675 0.7325  ;
        POLYGON 1.5625 0.625 1.9725 0.625 1.9725 0.69 1.5625 0.69  ;
    END
  END EN
  OBS
      LAYER metal1 ;
        POLYGON 0.7675 0.5175 1.3675 0.5175 1.3675 0.5825 0.7675 0.5825  ;
        POLYGON 0.9825 1.1125 1.2525 1.1125 1.2525 1.1525 1.6425 1.1525 1.6425 0.7575 1.8225 0.7575 1.8225 0.8225 1.7075 0.8225 1.7075 1.2175 1.1925 1.2175 1.1925 1.1775 0.9425 1.1775 0.9425 1.2025 0.9275 1.2025 0.9275 1.225 0.4275 1.225 0.4275 0.7 0.1175 0.7 0.1175 1.115 0.1225 1.115 0.1225 1.25 0.0525 1.25 0.0525 0.6525 0.0725 0.6525 0.0725 0.2675 0.1375 0.2675 0.1375 0.635 0.4925 0.635 0.4925 1.16 0.8775 1.16 0.8775 1.1175 0.9175 1.1175 0.9175 0.7975 1.0525 0.7975 1.0525 0.8625 0.9825 0.8625  ;
        POLYGON 2.0125 1.1075 2.0375 1.1075 2.0375 0.4925 1.5625 0.4925 1.5625 0.4275 2.0325 0.4275 2.0325 0.2675 2.0975 0.2675 2.0975 0.4675 2.1025 0.4675 2.1025 1.2425 2.0125 1.2425  ;
  END
END TBUF_X8

MACRO TINV_X1
  CLASS core ;
  FOREIGN TINV_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 0.76 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.235 1.315 0.235 0.92 0.3 0.92 0.3 1.315 0.76 1.315 0.76 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 0.76 -0.085 0.76 0.085 0.32 0.085 0.32 0.2925 0.255 0.2925 0.255 0.085 0 0.085  ;
    END
  END VSS
  PIN I
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.335 0.5375 0.4 0.5375 0.4 0.5975 0.5425 0.5975 0.5425 0.6725 0.335 0.6725  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 1.0175 0.63 1.0175 0.63 0.2125 0.695 0.2125 0.695 1.0825 0.4075 1.0825  ;
    END
  END ZN
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.18 0.6675 0.245 0.6675 0.245 0.7375 0.565 0.7375 0.565 0.8725 0.5 0.8725 0.5 0.8025 0.18 0.8025  ;
    END
  END EN
  OBS
      LAYER metal1 ;
        POLYGON 0.05 0.2125 0.115 0.2125 0.115 0.4075 0.5 0.4075 0.5 0.3375 0.565 0.3375 0.565 0.4725 0.115 0.4725 0.115 0.995 0.05 0.995  ;
  END
END TINV_X1

MACRO TLAT_X1
  CLASS core ;
  FOREIGN TLAT_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 2.66 BY 1.4 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.23 1.315 0.23 1.0425 0.295 1.0425 0.295 1.315 0.595 1.315 0.595 1.0675 0.66 1.0675 0.66 1.315 1.315 1.315 1.315 1.1025 1.45 1.1025 1.45 1.315 1.97 1.315 1.97 0.8725 2.035 0.8725 2.035 1.315 2.66 1.315 2.66 1.485 0 1.485  ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 2.3425 0.5625 2.365 0.5625 2.365 0.3675 2.43 0.3675 2.43 1.025 2.365 1.025 2.365 0.6975 2.3425 0.6975  ;
    END
  END Q
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 2.66 -0.085 2.66 0.085 2.055 0.085 2.055 0.4475 1.99 0.4475 1.99 0.085 1.43 0.085 1.43 0.175 1.295 0.175 1.295 0.085 0.64 0.085 0.64 0.21 0.575 0.21 0.575 0.085 0.33 0.085 0.33 0.3 0.195 0.3 0.195 0.085 0 0.085  ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.6325 0.5625 0.64 0.5625 0.64 0.34 0.78 0.34 0.78 0.405 0.705 0.405 0.705 0.74 0.775 0.74 0.775 0.805 0.64 0.805 0.64 0.6975 0.6325 0.6975  ;
    END
  END D
  PIN OE
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 1.3925 0.8375 1.55 0.8375 1.55 0.9025 1.4575 0.9025 1.4575 0.9775 1.3925 0.9775  ;
    END
  END OE
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.175 0.8075 0.3175 0.8075 0.3175 0.9775 0.2525 0.9775 0.2525 0.8725 0.175 0.8725  ;
    END
  END G
  OBS
      LAYER metal1 ;
        POLYGON 0.045 0.305 0.11 0.305 0.11 0.43 0.34 0.43 0.34 0.565 0.11 0.565 0.11 1.1725 0.045 1.1725  ;
        POLYGON 0.505 0.87 0.865 0.87 0.865 0.8325 1.115 0.8325 1.115 0.915 0.9125 0.915 0.9125 0.9225 0.905 0.9225 0.905 0.935 0.505 0.935 0.505 1.1725 0.44 1.1725 0.44 0.5125 0.42 0.5125 0.42 0.29 0.485 0.29 0.485 0.465 0.575 0.465 0.575 0.53 0.505 0.53  ;
        POLYGON 0.94 0.99 1.18 0.99 1.18 0.6375 1.14 0.6375 1.14 0.28 0.92 0.28 0.92 0.215 1.205 0.215 1.205 0.5775 1.215 0.5775 1.215 0.5825 1.645 0.5825 1.645 0.7175 1.245 0.7175 1.245 1.055 1.075 1.055 1.075 1.195 0.94 1.195  ;
        POLYGON 1.27 0.4525 1.795 0.4525 1.795 0.5175 1.775 0.5175 1.775 1.0025 1.71 1.0025 1.71 0.5175 1.27 0.5175  ;
        POLYGON 1.52 1.1825 1.84 1.1825 1.84 0.76 1.86 0.76 1.86 0.245 1.585 0.245 1.585 0.2225 1.5 0.2225 1.5 0.1575 1.635 0.1575 1.635 0.18 1.925 0.18 1.925 0.7425 2.26 0.7425 2.26 0.7475 2.3 0.7475 2.3 0.8825 2.235 0.8825 2.235 0.8075 1.905 0.8075 1.905 1.2475 1.52 1.2475  ;
  END
END TLAT_X1

MACRO XNOR2_X1
  CLASS core ;
  FOREIGN XNOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.2175 0.4575 0.76 0.4575 0.76 0.5925 0.2175 0.5925  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.085 1.315 0.085 1.175 0.15 1.175 0.15 1.315 0.46 1.315 0.46 1.175 0.525 1.175 0.525 1.315 1.03 1.315 1.03 1.175 1.095 1.175 1.095 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.525 0.085 0.525 0.3925 0.46 0.3925 0.46 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.4075 0.915 0.885 0.915 0.885 0.845 0.95 0.845 0.95 0.98 0.5425 0.98 0.5425 1.0825 0.4075 1.0825  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.655 1.115 0.8575 1.115 0.8575 1.045 1.015 1.045 1.015 0.5225 0.845 0.5225 0.845 0.3125 0.91 0.3125 0.91 0.4575 1.08 0.4575 1.08 1.11 0.9225 1.11 0.9225 1.2225 0.72 1.2225 0.72 1.25 0.655 1.25  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.655 0.1825 1.095 0.1825 1.095 0.3925 1.03 0.3925 1.03 0.2475 0.72 0.2475 0.72 0.3925 0.655 0.3925  ;
        POLYGON 0.085 0.3125 0.15 0.3125 0.15 0.715 0.61 0.715 0.61 0.85 0.545 0.85 0.545 0.78 0.335 0.78 0.335 1.25 0.27 1.25 0.27 0.78 0.1 0.78 0.1 0.7575 0.085 0.7575  ;
  END
END XNOR2_X1

MACRO XNOR2_X2
  CLASS core ;
  FOREIGN XNOR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.19 0.5025 0.2175 0.5025 0.2175 0.4575 0.3525 0.4575 0.3525 0.5725 0.745 0.5725 0.745 0.7075 0.68 0.7075 0.68 0.6375 0.19 0.6375  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.045 1.315 0.045 1.1875 0.11 1.1875 0.11 1.315 0.44 1.315 0.44 1.0475 0.505 1.0475 0.505 1.315 1.02 1.315 1.02 1.1875 1.085 1.1875 1.085 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 0.505 0.085 0.505 0.5075 0.44 0.5075 0.44 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.34 0.7025 0.405 0.7025 0.405 0.7725 0.875 0.7725 0.875 0.7425 0.94 0.7425 0.94 0.8775 0.9225 0.8775 0.9225 0.9425 0.7875 0.9425 0.7875 0.8375 0.34 0.8375  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.61 1.015 1.005 1.015 1.005 0.6375 0.905 0.6375 0.905 0.6325 0.865 0.6325 0.865 0.5225 0.7875 0.5225 0.7875 0.4575 0.795 0.4575 0.795 0.3125 0.93 0.3125 0.93 0.3775 0.86 0.3775 0.86 0.4525 0.93 0.4525 0.93 0.5725 1.07 0.5725 1.07 1.08 0.745 1.08 0.745 1.22 0.61 1.22  ;
    END
  END ZN
  OBS
      LAYER metal1 ;
        POLYGON 0.645 0.1825 1.085 0.1825 1.085 0.5075 1.02 0.5075 1.02 0.2475 0.71 0.2475 0.71 0.5075 0.645 0.5075  ;
        POLYGON 0.195 1.1625 0.265 1.1625 0.265 0.9675 0.045 0.9675 0.045 0.2875 0.11 0.2875 0.11 0.9025 0.565 0.9025 0.565 0.9675 0.33 0.9675 0.33 1.2275 0.195 1.2275  ;
  END
END XNOR2_X2

MACRO XOR2_X1
  CLASS core ;
  FOREIGN XOR2_X1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.805 0.8775 0.975 0.8775 0.975 0.3825 0.6575 0.3825 0.6575 0.3375 0.615 0.3375 0.615 0.1725 0.68 0.1725 0.68 0.2725 0.7225 0.2725 0.7225 0.3175 1.04 0.3175 1.04 0.9425 0.87 0.9425 0.87 1.02 0.805 1.02  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.19 0.76 0.72 0.76 0.72 0.9425 0.19 0.9425  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.42 1.315 0.42 1.0075 0.485 1.0075 0.485 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 1.055 0.085 1.055 0.2525 0.99 0.2525 0.99 0.085 0.485 0.085 0.485 0.2925 0.42 0.2925 0.42 0.085 0.11 0.085 0.11 0.2925 0.045 0.2925 0.045 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.305 0.5975 0.91 0.5975 0.91 0.765 0.845 0.765 0.845 0.6625 0.305 0.6625  ;
    END
  END B
  OBS
      LAYER metal1 ;
        POLYGON 0.615 1.0075 0.68 1.0075 0.68 1.085 0.99 1.085 0.99 1.0075 1.055 1.0075 1.055 1.15 0.615 1.15  ;
        POLYGON 0.045 0.43 0.23 0.43 0.23 0.1725 0.295 0.1725 0.295 0.43 0.505 0.43 0.505 0.395 0.57 0.395 0.57 0.43 0.57 0.495 0.57 0.53 0.505 0.53 0.505 0.495 0.11 0.495 0.11 1.02 0.045 1.02  ;
  END
END XOR2_X1

MACRO XOR2_X2
  CLASS core ;
  FOREIGN XOR2_X2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE NCSU_FreePDK_45nm ;
  SIZE 1.14 BY 1.4 ;
  PIN Z
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.7875 0.91 0.875 0.91 0.875 0.84 0.9925 0.84 0.9925 0.425 0.6325 0.425 0.6325 0.15 0.6975 0.15 0.6975 0.36 1.0575 0.36 1.0575 0.905 0.94 0.905 0.94 0.955 0.9225 0.955 0.9225 1.115 0.7875 1.115  ;
    END
  END Z
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.1925 0.78 0.81 0.78 0.81 0.845 0.5425 0.845 0.5425 0.9425 0.4075 0.9425 0.4075 0.915 0.1925 0.915  ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 1.315 0.4425 1.315 0.4425 1.05 0.5075 1.05 0.5075 1.315 1.14 1.315 1.14 1.485 0 1.485  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        POLYGON 0 -0.085 1.14 -0.085 1.14 0.085 1.0725 0.085 1.0725 0.285 1.0075 0.285 1.0075 0.085 0.4875 0.085 0.4875 0.375 0.4225 0.375 0.4225 0.085 0.1125 0.085 0.1125 0.375 0.0475 0.375 0.0475 0.085 0 0.085  ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        POLYGON 0.3425 0.58 0.4075 0.58 0.4075 0.65 0.8225 0.65 0.8225 0.5625 0.9275 0.5625 0.9275 0.715 0.3425 0.715  ;
    END
  END B
  OBS
      LAYER metal1 ;
        POLYGON 0.6325 0.97 0.6975 0.97 0.6975 1.18 1.0075 1.18 1.0075 0.97 1.0725 0.97 1.0725 1.245 0.6325 1.245  ;
        POLYGON 0.0475 0.495 0.0625 0.495 0.0625 0.4725 0.2325 0.4725 0.2325 0.255 0.2975 0.255 0.2975 0.45 0.5725 0.45 0.5725 0.585 0.5075 0.585 0.5075 0.515 0.2825 0.515 0.2825 0.5375 0.1125 0.5375 0.1125 1.2025 0.0475 1.2025  ;
  END
END XOR2_X2

END LIBRARY
#
# End of file
#
